library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
use WORK.constants.all;

entity TB_DRAM is
end TB_DRAM;

architecture TEST of TB_DRAM is
  constant NBITADDRESS : integer := NumBitMemoryAddress;
  constant NBITDATA : integer := NumBitMemoryWord;
  signal tb_address : std_logic_vector(NBITADDRESS-1 downto 0);
  signal tb_data_in : std_logic_vector(NBITDATA-1 downto 0);
  signal tb_write_enable : std_logic := '1';
  signal tb_read_enable : std_logic := '1';
  signal tb_data_out : std_logic_vector(NBITDATA-1 downto 0);

  component DRAM
  generic(MBIT : integer := NumBitMemoryWord;
          NBIT : integer := NumBitMemoryAddress);
  port(address : IN std_logic_vector(NBIT-1 downto 0);
       data_in : IN std_logic_vector(MBIT-1 downto 0);
       write_enable : IN std_logic;
       read_enable : IN std_logic;
       data_out : OUT std_logic_vector(MBIT-1 downto 0));
  end component;

  begin
    DUT : DRAM
    generic map(NBITDATA,NBITADDRESS)
    port map(tb_address,tb_data_in,tb_write_enable,tb_read_enable,tb_data_out);

    tb_data_in <= "11111111111111111111111111111111", "00000000000000000000000000000000" after 20 ns, "11111111111111111111111111111111" after 25 ns;
    tb_address <= "00000000";
    tb_write_enable <= '1','0' after 13 ns, '1' after 20 ns;
    tb_read_enable <= '0' after 4 ns, '1' after 13 ns,'0' after 20 ns, '1' after 25 ns;

  end TEST;

configuration CFG_TB_DRAM of TB_DRAM is
  for TEST
    for DUT : DRAM
      use configuration WORK.CFG_DRAM;
    end for;
  end for;
end CFG_TB_DRAM;
