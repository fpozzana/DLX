
module CU_HARDWIRED ( MUXA_CONTROL, MUXB_CONTROL, ALU_OPCODE, DRAM_WE, DRAM_RE, 
        WB_MUX_SEL, JAL_SEL, RF_WE, OPCODE, FUNC, Clk, Rst );
  output [3:0] ALU_OPCODE;
  input [5:0] OPCODE;
  input [10:0] FUNC;
  input Clk, Rst;
  output MUXA_CONTROL, MUXB_CONTROL, DRAM_WE, DRAM_RE, WB_MUX_SEL, JAL_SEL,
         RF_WE;

  assign MUXA_CONTROL = 1'b0;
  assign MUXB_CONTROL = 1'b0;
  assign ALU_OPCODE[3] = 1'b0;
  assign ALU_OPCODE[2] = 1'b0;
  assign ALU_OPCODE[1] = 1'b0;
  assign ALU_OPCODE[0] = 1'b0;
  assign DRAM_WE = 1'b0;
  assign DRAM_RE = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign JAL_SEL = 1'b0;
  assign RF_WE = 1'b0;

endmodule


module FD_0 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_302 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_301 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_300 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_299 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_298 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_297 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_296 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_295 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_294 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_293 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_292 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_291 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_290 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_289 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_288 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_287 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_286 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_285 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_284 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_283 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_282 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_281 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_280 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_279 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_278 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_277 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_276 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_275 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_274 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_273 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_272 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_0 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n18, n19, n20;

  FD_0 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n20), .Q(Q[0]) );
  FD_302 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n18), .Q(Q[1]) );
  FD_301 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n18), .Q(Q[2]) );
  FD_300 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n18), .Q(Q[3]) );
  FD_299 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n18), .Q(Q[4]) );
  FD_298 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n18), .Q(Q[5]) );
  FD_297 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n18), .Q(Q[6]) );
  FD_296 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n18), .Q(Q[7]) );
  FD_295 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n18), .Q(Q[8]) );
  FD_294 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n18), .Q(Q[9]) );
  FD_293 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n18), .Q(Q[10]) );
  FD_292 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n18), .Q(Q[11]) );
  FD_291 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n18), .Q(Q[12]) );
  FD_290 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n19), .Q(Q[13]) );
  FD_289 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n19), .Q(Q[14]) );
  FD_288 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n19), .Q(Q[15]) );
  FD_287 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n19), .Q(Q[16]) );
  FD_286 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n19), .Q(Q[17]) );
  FD_285 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n19), .Q(Q[18]) );
  FD_284 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n19), .Q(Q[19]) );
  FD_283 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n19), .Q(Q[20]) );
  FD_282 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n19), .Q(Q[21]) );
  FD_281 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n19), .Q(Q[22]) );
  FD_280 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n19), .Q(Q[23]) );
  FD_279 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n19), .Q(Q[24]) );
  FD_278 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n20), .Q(Q[25]) );
  FD_277 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n20), .Q(Q[26]) );
  FD_276 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n20), .Q(Q[27]) );
  FD_275 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n20), .Q(Q[28]) );
  FD_274 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n20), .Q(Q[29]) );
  FD_273 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n20), .Q(Q[30]) );
  FD_272 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n20), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n18) );
  BUF_X1 U2 ( .A(RESET), .Z(n19) );
  BUF_X1 U3 ( .A(RESET), .Z(n20) );
endmodule


module FD_271 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_270 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_269 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_268 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_267 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_266 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_265 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_264 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_263 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_262 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_261 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_260 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_259 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_258 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_257 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_256 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_255 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_254 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_253 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_252 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_251 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_250 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_249 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_248 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_247 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_246 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n8;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n8), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n8) );
endmodule


module FD_245 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_244 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_243 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_242 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_241 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_240 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_8 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_271 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_270 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_269 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_268 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_267 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_266 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_265 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_264 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_263 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_262 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_261 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_260 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_259 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_258 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_257 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_256 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_255 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_254 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_253 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_252 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_251 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_250 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_249 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_248 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_247 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_246 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_245 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_244 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_243 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_242 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_241 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_240 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FETCH_STAGE_numbit32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n4, n6, n7, n8, n10, n13, n16, n17, n18, n19,
         n20, n23, n25, n27, n30, n31, n32, n34, n35, n36, n37, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n57,
         n61, n66, n69, n70, n71, n72, n75, n77, n79, n80, n82, n85, n88, n91,
         n94, n95, n96, n97, n98, n99, n101, n104, n106, n107, n110, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND3_X1 U25 ( .A1(A[19]), .A2(A[18]), .A3(n10), .ZN(n13) );
  NAND3_X1 U36 ( .A1(A[6]), .A2(n61), .A3(n107), .ZN(n23) );
  NAND3_X1 U55 ( .A1(A[23]), .A2(A[22]), .A3(n32), .ZN(n35) );
  NAND3_X1 U56 ( .A1(A[19]), .A2(A[18]), .A3(n10), .ZN(n72) );
  XOR2_X1 U58 ( .A(n37), .B(A[23]), .Z(SUM[23]) );
  NAND3_X1 U64 ( .A1(A[10]), .A2(n25), .A3(A[11]), .ZN(n96) );
  NAND3_X1 U67 ( .A1(A[23]), .A2(A[22]), .A3(n32), .ZN(n71) );
  XOR2_X1 U73 ( .A(A[14]), .B(n101), .Z(SUM[14]) );
  XOR2_X1 U74 ( .A(n55), .B(n177), .Z(SUM[7]) );
  XOR2_X1 U75 ( .A(A[5]), .B(n52), .Z(SUM[5]) );
  XOR2_X1 U76 ( .A(n91), .B(A[18]), .Z(SUM[18]) );
  XOR2_X1 U77 ( .A(A[2]), .B(A[3]), .Z(SUM[3]) );
  XOR2_X1 U85 ( .A(n44), .B(n188), .Z(SUM[12]) );
  XOR2_X1 U86 ( .A(A[8]), .B(n50), .Z(SUM[8]) );
  XOR2_X1 U87 ( .A(n45), .B(n181), .Z(SUM[13]) );
  XOR2_X1 U88 ( .A(n104), .B(n179), .Z(SUM[11]) );
  XOR2_X1 U89 ( .A(n31), .B(n187), .Z(SUM[16]) );
  XOR2_X1 U90 ( .A(n106), .B(A[10]), .Z(SUM[10]) );
  XOR2_X1 U91 ( .A(n53), .B(n180), .Z(SUM[9]) );
  XOR2_X1 U102 ( .A(n2), .B(A[26]), .Z(SUM[26]) );
  XOR2_X1 U103 ( .A(n51), .B(A[17]), .Z(SUM[17]) );
  NAND3_X1 U132 ( .A1(A[13]), .A2(A[12]), .A3(A[14]), .ZN(n97) );
  NAND3_X1 U133 ( .A1(A[5]), .A2(A[7]), .A3(A[4]), .ZN(n98) );
  XOR2_X1 U2 ( .A(n110), .B(A[29]), .Z(SUM[29]) );
  NAND3_X1 U7 ( .A1(A[30]), .A2(A[29]), .A3(n8), .ZN(n34) );
  XOR2_X1 U8 ( .A(A[4]), .B(n61), .Z(SUM[4]) );
  XOR2_X1 U9 ( .A(n39), .B(A[15]), .Z(SUM[15]) );
  AND2_X1 U3 ( .A1(n69), .A2(n42), .ZN(n43) );
  XNOR2_X1 U4 ( .A(n1), .B(n185), .ZN(SUM[24]) );
  AND2_X1 U5 ( .A1(n82), .A2(n49), .ZN(n1) );
  NAND2_X1 U6 ( .A1(n88), .A2(n6), .ZN(n40) );
  NOR2_X1 U10 ( .A1(n31), .A2(n182), .ZN(n6) );
  NOR2_X1 U11 ( .A1(n79), .A2(n47), .ZN(n46) );
  NAND2_X1 U12 ( .A1(n7), .A2(n88), .ZN(n48) );
  NOR2_X1 U13 ( .A1(n31), .A2(n182), .ZN(n7) );
  NAND2_X1 U14 ( .A1(n82), .A2(n49), .ZN(n79) );
  AND2_X1 U15 ( .A1(n70), .A2(n49), .ZN(n42) );
  OR2_X1 U16 ( .A1(n186), .A2(n183), .ZN(n41) );
  XNOR2_X1 U17 ( .A(n85), .B(n186), .ZN(SUM[22]) );
  NOR2_X1 U18 ( .A1(n48), .A2(n183), .ZN(n85) );
  OR2_X1 U19 ( .A1(n44), .A2(n188), .ZN(n45) );
  AND2_X1 U20 ( .A1(n95), .A2(n17), .ZN(n49) );
  NAND2_X1 U21 ( .A1(n95), .A2(n17), .ZN(n31) );
  AND2_X1 U22 ( .A1(n30), .A2(n17), .ZN(n51) );
  NOR2_X1 U23 ( .A1(n44), .A2(n20), .ZN(n101) );
  OR2_X1 U24 ( .A1(n188), .A2(n181), .ZN(n20) );
  XNOR2_X1 U26 ( .A(A[30]), .B(n66), .ZN(SUM[30]) );
  NAND2_X1 U27 ( .A1(n43), .A2(A[29]), .ZN(n66) );
  AND2_X1 U28 ( .A1(n69), .A2(n42), .ZN(n110) );
  XNOR2_X1 U29 ( .A(A[31]), .B(n34), .ZN(SUM[31]) );
  AND4_X1 U30 ( .A1(A[27]), .A2(A[25]), .A3(A[26]), .A4(A[24]), .ZN(n16) );
  AND2_X1 U31 ( .A1(A[28]), .A2(n16), .ZN(n69) );
  AND4_X1 U32 ( .A1(A[28]), .A2(n70), .A3(n16), .A4(n49), .ZN(n8) );
  XNOR2_X1 U33 ( .A(n77), .B(A[27]), .ZN(SUM[27]) );
  NAND2_X1 U34 ( .A1(n46), .A2(A[26]), .ZN(n77) );
  NOR2_X1 U35 ( .A1(n71), .A2(n72), .ZN(n82) );
  NOR2_X1 U37 ( .A1(n35), .A2(n13), .ZN(n70) );
  NOR2_X1 U38 ( .A1(n40), .A2(n41), .ZN(n37) );
  NOR2_X1 U39 ( .A1(n79), .A2(n47), .ZN(n2) );
  INV_X1 U40 ( .A(A[20]), .ZN(n182) );
  INV_X1 U41 ( .A(A[24]), .ZN(n185) );
  INV_X1 U42 ( .A(A[22]), .ZN(n186) );
  INV_X1 U43 ( .A(A[21]), .ZN(n183) );
  AND2_X1 U44 ( .A1(A[21]), .A2(A[20]), .ZN(n32) );
  OR2_X1 U45 ( .A1(n184), .A2(n185), .ZN(n47) );
  INV_X1 U46 ( .A(A[25]), .ZN(n184) );
  XNOR2_X1 U47 ( .A(n80), .B(A[25]), .ZN(SUM[25]) );
  NAND2_X1 U48 ( .A1(n1), .A2(A[24]), .ZN(n80) );
  XNOR2_X1 U49 ( .A(n48), .B(A[21]), .ZN(SUM[21]) );
  XNOR2_X1 U50 ( .A(n75), .B(A[28]), .ZN(SUM[28]) );
  NAND2_X1 U51 ( .A1(n1), .A2(n16), .ZN(n75) );
  AND2_X1 U52 ( .A1(A[8]), .A2(A[9]), .ZN(n25) );
  XNOR2_X1 U53 ( .A(n36), .B(A[19]), .ZN(SUM[19]) );
  NAND2_X1 U54 ( .A1(n51), .A2(n27), .ZN(n36) );
  AND3_X1 U57 ( .A1(A[19]), .A2(A[18]), .A3(n10), .ZN(n88) );
  NOR2_X1 U59 ( .A1(n96), .A2(n97), .ZN(n95) );
  NOR2_X1 U60 ( .A1(n53), .A2(n180), .ZN(n106) );
  INV_X1 U61 ( .A(A[11]), .ZN(n179) );
  AND2_X1 U62 ( .A1(A[14]), .A2(n101), .ZN(n39) );
  AND2_X1 U63 ( .A1(n30), .A2(n19), .ZN(n91) );
  AND2_X1 U65 ( .A1(n94), .A2(A[15]), .ZN(n17) );
  NOR2_X1 U66 ( .A1(n98), .A2(n99), .ZN(n94) );
  NAND2_X1 U68 ( .A1(A[6]), .A2(n61), .ZN(n99) );
  OR2_X1 U69 ( .A1(n23), .A2(n96), .ZN(n44) );
  INV_X1 U70 ( .A(A[9]), .ZN(n180) );
  INV_X1 U71 ( .A(A[12]), .ZN(n188) );
  AND2_X1 U72 ( .A1(A[17]), .A2(A[16]), .ZN(n10) );
  INV_X1 U78 ( .A(A[13]), .ZN(n181) );
  OR2_X1 U79 ( .A1(n53), .A2(n4), .ZN(n104) );
  NAND2_X1 U80 ( .A1(A[10]), .A2(A[9]), .ZN(n4) );
  AND2_X1 U81 ( .A1(n95), .A2(A[16]), .ZN(n30) );
  AND2_X1 U82 ( .A1(A[18]), .A2(A[17]), .ZN(n27) );
  INV_X1 U83 ( .A(A[16]), .ZN(n187) );
  XNOR2_X1 U84 ( .A(n18), .B(A[20]), .ZN(SUM[20]) );
  NAND2_X1 U92 ( .A1(n88), .A2(n49), .ZN(n18) );
  AND2_X1 U93 ( .A1(n17), .A2(A[17]), .ZN(n19) );
  NAND2_X1 U94 ( .A1(A[6]), .A2(n57), .ZN(n55) );
  AND2_X1 U95 ( .A1(A[3]), .A2(A[2]), .ZN(n61) );
  NAND2_X1 U96 ( .A1(n50), .A2(A[8]), .ZN(n53) );
  AND2_X1 U97 ( .A1(n52), .A2(A[5]), .ZN(n57) );
  AND3_X1 U98 ( .A1(A[6]), .A2(n61), .A3(n107), .ZN(n50) );
  XNOR2_X1 U99 ( .A(n178), .B(n57), .ZN(SUM[6]) );
  INV_X1 U100 ( .A(A[6]), .ZN(n178) );
  AND3_X1 U101 ( .A1(A[7]), .A2(A[5]), .A3(A[4]), .ZN(n107) );
  AND2_X1 U104 ( .A1(n61), .A2(A[4]), .ZN(n52) );
  INV_X1 U105 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U106 ( .A(A[7]), .ZN(n177) );
endmodule


module FETCH_STAGE_numbit32 ( program_counter, to_IR, clk, reset, to_IRAM, 
        npc_out, instruction_reg_out, instruction_fetched );
  input [31:0] program_counter;
  input [31:0] to_IR;
  output [31:0] to_IRAM;
  output [31:0] npc_out;
  output [31:0] instruction_reg_out;
  output [31:0] instruction_fetched;
  input clk, reset;
  wire   N0, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n47, n48, n49
;
  wire   [31:0] adder_out;
  assign to_IRAM[31] = 1'b0;
  assign to_IRAM[30] = 1'b0;
  assign instruction_fetched[31] = to_IR[31];
  assign instruction_fetched[30] = to_IR[30];
  assign instruction_fetched[29] = to_IR[29];
  assign instruction_fetched[28] = to_IR[28];
  assign instruction_fetched[27] = to_IR[27];
  assign instruction_fetched[26] = to_IR[26];
  assign instruction_fetched[25] = to_IR[25];
  assign instruction_fetched[24] = to_IR[24];
  assign instruction_fetched[23] = to_IR[23];
  assign instruction_fetched[22] = to_IR[22];
  assign instruction_fetched[21] = to_IR[21];
  assign instruction_fetched[20] = to_IR[20];
  assign instruction_fetched[19] = to_IR[19];
  assign instruction_fetched[18] = to_IR[18];
  assign instruction_fetched[17] = to_IR[17];
  assign instruction_fetched[16] = to_IR[16];
  assign instruction_fetched[15] = to_IR[15];
  assign instruction_fetched[14] = to_IR[14];
  assign instruction_fetched[13] = to_IR[13];
  assign instruction_fetched[12] = to_IR[12];
  assign instruction_fetched[11] = to_IR[11];
  assign instruction_fetched[10] = to_IR[10];
  assign instruction_fetched[9] = to_IR[9];
  assign instruction_fetched[8] = to_IR[8];
  assign instruction_fetched[7] = to_IR[7];
  assign instruction_fetched[6] = to_IR[6];
  assign instruction_fetched[5] = to_IR[5];
  assign instruction_fetched[4] = to_IR[4];
  assign instruction_fetched[3] = to_IR[3];
  assign instruction_fetched[2] = to_IR[2];
  assign instruction_fetched[1] = to_IR[1];
  assign instruction_fetched[0] = to_IR[0];

  DLH_X1 \to_IRAM_reg[29]  ( .G(n47), .D(program_counter[31]), .Q(to_IRAM[29])
         );
  DLH_X1 \to_IRAM_reg[28]  ( .G(n47), .D(program_counter[30]), .Q(to_IRAM[28])
         );
  DLH_X1 \to_IRAM_reg[27]  ( .G(n47), .D(program_counter[29]), .Q(to_IRAM[27])
         );
  DLH_X1 \to_IRAM_reg[26]  ( .G(n48), .D(program_counter[28]), .Q(to_IRAM[26])
         );
  DLH_X1 \to_IRAM_reg[25]  ( .G(n48), .D(program_counter[27]), .Q(to_IRAM[25])
         );
  DLH_X1 \to_IRAM_reg[24]  ( .G(n48), .D(program_counter[26]), .Q(to_IRAM[24])
         );
  DLH_X1 \to_IRAM_reg[23]  ( .G(n48), .D(program_counter[25]), .Q(to_IRAM[23])
         );
  DLH_X1 \to_IRAM_reg[22]  ( .G(n48), .D(program_counter[24]), .Q(to_IRAM[22])
         );
  DLH_X1 \to_IRAM_reg[21]  ( .G(n48), .D(program_counter[23]), .Q(to_IRAM[21])
         );
  DLH_X1 \to_IRAM_reg[20]  ( .G(n48), .D(program_counter[22]), .Q(to_IRAM[20])
         );
  DLH_X1 \to_IRAM_reg[19]  ( .G(n48), .D(program_counter[21]), .Q(to_IRAM[19])
         );
  DLH_X1 \to_IRAM_reg[18]  ( .G(n49), .D(program_counter[20]), .Q(to_IRAM[18])
         );
  DLH_X1 \to_IRAM_reg[17]  ( .G(n49), .D(program_counter[19]), .Q(to_IRAM[17])
         );
  DLH_X1 \to_IRAM_reg[16]  ( .G(n49), .D(program_counter[18]), .Q(to_IRAM[16])
         );
  DLH_X1 \to_IRAM_reg[15]  ( .G(n49), .D(program_counter[17]), .Q(to_IRAM[15])
         );
  DLH_X1 \to_IRAM_reg[14]  ( .G(n49), .D(program_counter[16]), .Q(to_IRAM[14])
         );
  DLH_X1 \to_IRAM_reg[13]  ( .G(n48), .D(program_counter[15]), .Q(to_IRAM[13])
         );
  DLH_X1 \to_IRAM_reg[12]  ( .G(n48), .D(program_counter[14]), .Q(to_IRAM[12])
         );
  DLH_X1 \to_IRAM_reg[11]  ( .G(n48), .D(program_counter[13]), .Q(to_IRAM[11])
         );
  DLH_X1 \to_IRAM_reg[10]  ( .G(n47), .D(program_counter[12]), .Q(to_IRAM[10])
         );
  DLH_X1 \to_IRAM_reg[9]  ( .G(n47), .D(program_counter[11]), .Q(to_IRAM[9])
         );
  DLH_X1 \to_IRAM_reg[8]  ( .G(n47), .D(program_counter[10]), .Q(to_IRAM[8])
         );
  DLH_X1 \to_IRAM_reg[7]  ( .G(n47), .D(program_counter[9]), .Q(to_IRAM[7]) );
  DLH_X1 \to_IRAM_reg[6]  ( .G(n47), .D(program_counter[8]), .Q(to_IRAM[6]) );
  DLH_X1 \to_IRAM_reg[5]  ( .G(n47), .D(program_counter[7]), .Q(to_IRAM[5]) );
  DLH_X1 \to_IRAM_reg[4]  ( .G(n47), .D(program_counter[6]), .Q(to_IRAM[4]) );
  DLH_X1 \to_IRAM_reg[3]  ( .G(n47), .D(program_counter[5]), .Q(to_IRAM[3]) );
  DLH_X1 \to_IRAM_reg[2]  ( .G(n49), .D(program_counter[4]), .Q(to_IRAM[2]) );
  DLH_X1 \to_IRAM_reg[1]  ( .G(n49), .D(program_counter[3]), .Q(to_IRAM[1]) );
  DLH_X1 \to_IRAM_reg[0]  ( .G(n49), .D(program_counter[2]), .Q(to_IRAM[0]) );
  REGISTER_GENERIC_NBIT32_0 NPC ( .D(adder_out), .CK(clk), .RESET(reset), .Q(
        npc_out) );
  REGISTER_GENERIC_NBIT32_8 IR ( .D(to_IR), .CK(clk), .RESET(reset), .Q(
        instruction_reg_out) );
  FETCH_STAGE_numbit32_DW01_add_2 add_51 ( .A(program_counter), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(adder_out) );
  BUF_X1 U5 ( .A(N0), .Z(n48) );
  BUF_X1 U7 ( .A(N0), .Z(n47) );
  BUF_X1 U8 ( .A(N0), .Z(n49) );
  NOR4_X1 U11 ( .A1(program_counter[21]), .A2(program_counter[20]), .A3(
        program_counter[19]), .A4(program_counter[18]), .ZN(n12) );
  NOR4_X1 U12 ( .A1(program_counter[9]), .A2(program_counter[8]), .A3(
        program_counter[7]), .A4(program_counter[31]), .ZN(n17) );
  NOR3_X1 U13 ( .A1(program_counter[15]), .A2(program_counter[17]), .A3(
        program_counter[16]), .ZN(n11) );
  NOR3_X1 U14 ( .A1(program_counter[28]), .A2(program_counter[30]), .A3(
        program_counter[29]), .ZN(n16) );
  NOR3_X1 U15 ( .A1(program_counter[25]), .A2(program_counter[27]), .A3(
        program_counter[26]), .ZN(n15) );
  NOR3_X1 U16 ( .A1(program_counter[12]), .A2(program_counter[14]), .A3(
        program_counter[13]), .ZN(n10) );
  NOR3_X1 U17 ( .A1(n13), .A2(program_counter[11]), .A3(program_counter[10]), 
        .ZN(n9) );
  AND4_X1 U18 ( .A1(program_counter[6]), .A2(program_counter[5]), .A3(
        program_counter[4]), .A4(program_counter[3]), .ZN(n13) );
  NOR2_X1 U19 ( .A1(n7), .A2(n8), .ZN(N0) );
  NAND4_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .ZN(n7) );
  NAND4_X1 U21 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n8) );
  NOR3_X1 U22 ( .A1(program_counter[22]), .A2(program_counter[24]), .A3(
        program_counter[23]), .ZN(n14) );
endmodule


module SIGN_EXTENTION ( D, Q );
  input [15:0] D;
  output [31:0] Q;
  wire   \Q[31] , \Q[19] ;
  assign Q[14] = D[14];
  assign Q[13] = D[13];
  assign Q[12] = D[12];
  assign Q[11] = D[11];
  assign Q[10] = D[10];
  assign Q[9] = D[9];
  assign Q[8] = D[8];
  assign Q[7] = D[7];
  assign Q[6] = D[6];
  assign Q[5] = D[5];
  assign Q[4] = D[4];
  assign Q[3] = D[3];
  assign Q[2] = D[2];
  assign Q[1] = D[1];
  assign Q[0] = D[0];
  assign Q[20] = \Q[31] ;
  assign Q[21] = \Q[31] ;
  assign Q[22] = \Q[31] ;
  assign Q[23] = \Q[31] ;
  assign Q[24] = \Q[31] ;
  assign Q[25] = \Q[31] ;
  assign Q[26] = \Q[31] ;
  assign Q[27] = \Q[31] ;
  assign Q[28] = \Q[31] ;
  assign Q[29] = \Q[31] ;
  assign Q[30] = \Q[31] ;
  assign Q[31] = \Q[31] ;
  assign Q[15] = \Q[19] ;
  assign Q[16] = \Q[19] ;
  assign Q[17] = \Q[19] ;
  assign Q[18] = \Q[19] ;
  assign Q[19] = \Q[19] ;

  BUF_X1 U1 ( .A(D[15]), .Z(\Q[31] ) );
  BUF_X1 U2 ( .A(D[15]), .Z(\Q[19] ) );
endmodule


module REGISTER_FILE_numBit_data32_numBit_address5_numBit_registers32 ( CK, 
        Reset, Write_enable, Write_address, Read_one_address, Read_two_address, 
        Data_in, Data_one_out, Data_two_out );
  input [4:0] Write_address;
  input [4:0] Read_one_address;
  input [4:0] Read_two_address;
  input [31:0] Data_in;
  output [31:0] Data_one_out;
  output [31:0] Data_two_out;
  input CK, Reset, Write_enable;
  wire   N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N993,
         N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         n1155, n1156, n1164, n1165, n1166, n1169, n1173, n1174, n1175, n1179,
         n1180, n1181, n1183, n1184, n1185, n1186, n1187, n1190, n1191, n1192,
         n1193, n1195, n1197, n1198, n1199, n1200, n1203, n1204, n1206, n1207,
         n1208, n1210, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1223, n1225, n1226, n1228, n1233, n1235, n1236, n1237, n1238, n1240,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251, n1253,
         n1254, n1256, n1259, n1261, n1262, n1263, n1264, n1266, n1267, n1270,
         n1271, n1273, n1283, n1293, n1294, n1303, n1315, n1318, n1320, n1323,
         n1325, n1326, n1327, n1328, n1330, n1331, n1335, n1337, n1343, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1383, n1385, n1386, n1388, n1389,
         n1390, n1391, n1394, n1396, n1399, n1400, n1401, n1402, n1404, n1405,
         n1406, n1407, n1408, n1409, n1411, n1419, n1421, n1422, n1430, n1431,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1450, n1451, n1452,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1635, n1636, n1637,
         n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1648, n1649,
         n1651, n1653, n1654, n1655, n1659, n1660, n1661, n1664, n1665, n1667,
         n1668, n1669, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1685, n1686, n1687, n1689, n1691, n1692, n1693, n1695,
         n1700, n1701, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1713,
         n1714, n1717, n1719, n1721, n1723, n1724, n1725, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1775, n1778, n1785, n1791, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1827, n1829, n1833, n1834,
         n1837, n1838, n1846, n1847, n1855, n1858, n1859, n1863, n1869, n1870,
         n1876, n1878, n1879, n1880, n1882, n1886, n1887, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1936, n1937, n1939, n1940, n1941, n1943, n1944, n1946,
         n1947, n1948, n1949, n1950, n1951, n1955, n1956, n1957, n1958, n1960,
         n1961, n1962, n1963, n1964, n1967, n1968, n1969, n1970, n1971, n1973,
         n1974, n1977, n1979, n1980, n1981, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2051, n2052, n2053, n2054, n2056, n2057, n2058, n2060,
         n2063, n2064, n2065, n2066, n2067, n2069, n2073, n2075, n2076, n2077,
         n2079, n2080, n2081, n2093, n2094, n2102, n2103, n2114, n2115, n2116,
         n2117, n2119, n2121, n2124, n2125, n2126, n2129, n2132, n2133, n2134,
         n2135, n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n7813, n7821, n7822, n7830, n7831, n8079, n8080, n8085, n8086, n8100,
         n3147, n3203, n3208, n3224, n3225, n3226, n3227, n3228, n3229, n3240,
         n3242, n3310, n3311, n3329, n3333, n3335, n3337, n3354, n3356, n3358,
         n3360, n3362, n3381, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9347, n9348, n9349, n9350, n9356, n9357, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9378, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9411, n9417, n9418, n9419, n9420, n9421, n9433, n9434, n9435, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9462, n9466, n9467, n9468, n9469, n9470, n9472,
         n9473, n9478, n9479, n9480, n9481, n9482, n9483, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9500, n9502, n9503, n9506, n9523, n9524,
         n9525, n9526, n9527, n9528, n9537, n9538, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9558, n9559, n9560,
         n9562, n9563, n9566, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9579, n9580, n9581, n9582, n9583, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9612, n9613, n9614, n9615, n9627, n9629, n9630, n9632, n9640,
         n9641, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9655, n9656, n9659, n9660, n9661, n9662, n9664, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9681, n9683, n9684, n9685,
         n9721, n9722, n9723, n9725, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9754, n9759, n9760, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9781, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9803, n9811, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9835, n9836, n9837, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9856, n9857, n9858, n9860, n9861, n9862, n9863, n9864, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9890, n9891, n3053, n3055,
         n3060, n3061, n3062, n3079, n3083, n3084, n3085, n3088, n3089, n3091,
         n3094, n3095, n3101, n3106, n3117, n3118, n3119, n3120, n3121, n3122,
         n3128, n3129, n3130, n3131, n3136, n3137, n3138, n3146, n3148, n3149,
         n3153, n3156, n3158, n3159, n3160, n3167, n3180, n3181, n3182, n3193,
         n3194, n3213, n3214, n3215, n3216, n3217, n3218, n3220, n3221, n3222,
         n3223, n3230, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3241, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3265, n3266, n3267, n3268, n3269, n3275, n3282, n3283,
         n3284, n3285, n3289, n3290, n3291, n3292, n3293, n3295, n3296, n3297,
         n3299, n3303, n3304, n3305, n3312, n3320, n3321, n3322, n3323, n3324,
         n3325, n3341, n3344, n3346, n3347, n3348, n3351, n3352, n3353, n3355,
         n3357, n3359, n3361, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3379, n3382, n3383, n3594,
         n3629, n3630, n3631, n3632, n3633, n3635, n3637, n3639, n3640, n3641,
         n3642, n3643, n3650, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3665, n3667, n3669, n3671, n3673, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3688, n3689, n3692, n3693, n3697, n3698, n3699,
         n3700, n3703, n3704, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3716, n3718, n3720, n3721, n3722, n3723, n3724, n3725,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3093,
         n3098, n3111, n3112, n3113, n3116, n3127, n3135, n3139, n3140, n3141,
         n3142, n3143, n3144, n3178, n3184, n3185, n3188, n3189, n3201, n3207,
         n3286, n3298, n3300, n3301, n3308, n3314, n3316, n3328, n3330, n3332,
         n3380, n3664, n3670, n3672, n3702, n3726, n3789, n3795, n3796, n3799,
         n3801, n3805, n3807, n3808, n3809, n3810, n3812, n3814, n3815, n3817,
         n3819, n3820, n3821, n3822, n3824, n3826, n3827, n3828, n3829, n3830,
         n3833, n3834, n3835, n3836, n3837, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3853, n3854, n3856, n3858,
         n3861, n3864, n3866, n3868, n3875, n3881, n3884, n3895, n3896, n3897,
         n3898, n3900, n3903, n3909, n3916, n3917, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1095, n1097,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1117, n1118, n1119, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1167, n1168, n1170, n1171, n1172, n1176, n1177, n1178, n1182, n1188,
         n1189, n1194, n1196, n1201, n1202, n1205, n1209, n1211, n1212, n1213,
         n1222, n1224, n1227, n1229, n1230, n1231, n1232, n1234, n1239, n1241,
         n1250, n1252, n1255, n1257, n1258, n1260, n1265, n1268, n1269, n1272,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1319,
         n1321, n1322, n1324, n1329, n1332, n1333, n1334, n1336, n1338, n1339,
         n1340, n1341, n1342, n1344, n1345, n1382, n1384, n1387, n1392, n1393,
         n1395, n1397, n1398, n1403, n1410, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1420, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1432, n1433, n1434, n1435, n1437, n1438, n1439, n1440, n1441, n1449,
         n1453, n1454, n1463, n1471, n1634, n1639, n1647, n1650, n1652, n1656,
         n1657, n1658, n1662, n1663, n1670, n1671, n1672, n1683, n1684, n1688,
         n1690, n1694, n1696, n1697, n1698, n1699, n1702, n1703, n1704, n1712,
         n1715, n1716, n1718, n1720, n1722, n1726, n1727, n1737, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1776, n1777, n1779, n1780, n1781, n1782, n1783, n1784, n1786,
         n1787, n1788, n1789, n1790, n1792, n1793, n1826, n1828, n1830, n1831,
         n1832, n1835, n1836, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1856, n1857, n1860,
         n1861, n1862, n1864, n1865, n1866, n1867, n1868, n1871, n1872, n1873,
         n1874, n1875, n1877, n1881, n1883, n1884, n1885, n1888, n1889, n1935,
         n1938, n1942, n1945, n1952, n1953, n1954, n1959, n1965, n1966, n1972,
         n1975, n1976, n1978, n1982, n2050, n2055, n2059, n2061, n2062, n2068,
         n2070, n2071, n2072, n2074, n2078, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2118, n2120, n2122, n2123, n2127, n2128, n2130,
         n2131, n2137, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3054,
         n3056, n3057, n3058, n3059, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3080, n3081, n3082, n3086, n3087, n3092,
         n3099, n3100, n3102, n3103, n3104, n3105, n3107, n3108, n3109, n3110,
         n3114, n3115, n3123, n3124, n3125, n3126, n3132, n3133, n3134, n3150,
         n3151, n3152, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3176,
         n3177, n3186, n3187, n3191, n3192, n3196, n3202, n3209, n3211, n3212,
         n3219, n3231, n3264, n3271, n3272, n3273, n3276, n3277, n3278, n3279,
         n3280, n3281, n3287, n3288, n3302, n3306, n3307, n3309, n3313, n3315,
         n3317, n3319, n3331, n3339, n3340, n3343, n3345, n3349, n3378, n3628,
         n3634, n3638, n3644, n3645, n3649, n3659, n3660, n3663, n3666, n3684,
         n3685, n3696, n3790, n3818, n3831, n3832, n3839, n3851, n3855, n3865,
         n3867, n3869, n3873, n3876, n3877, n3880, n3883, n3886, n3888, n3889,
         n3891, n3892, n3894, n3899, n3914, n3918, n3919, n3920, n3921, n3922,
         n3924, n3925, n3939, n3941, n3943, n3944, n3946, n3947, n3948, n3951,
         n3952, n3953, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314;

  DLH_X1 \Data_one_out_reg[31]  ( .G(1'b1), .D(N991), .Q(Data_one_out[31]) );
  DLH_X1 \Data_one_out_reg[30]  ( .G(1'b1), .D(N990), .Q(Data_one_out[30]) );
  DLH_X1 \Data_one_out_reg[29]  ( .G(1'b1), .D(N989), .Q(Data_one_out[29]) );
  DLH_X1 \Data_one_out_reg[28]  ( .G(1'b1), .D(N988), .Q(Data_one_out[28]) );
  DLH_X1 \Data_one_out_reg[27]  ( .G(1'b1), .D(N987), .Q(Data_one_out[27]) );
  DLH_X1 \Data_one_out_reg[26]  ( .G(1'b1), .D(N986), .Q(Data_one_out[26]) );
  DLH_X1 \Data_one_out_reg[25]  ( .G(1'b1), .D(N985), .Q(Data_one_out[25]) );
  DLH_X1 \Data_one_out_reg[23]  ( .G(1'b1), .D(N983), .Q(Data_one_out[23]) );
  DLH_X1 \Data_one_out_reg[21]  ( .G(1'b1), .D(N981), .Q(Data_one_out[21]) );
  DLH_X1 \Data_one_out_reg[20]  ( .G(1'b1), .D(N980), .Q(Data_one_out[20]) );
  DLH_X1 \Data_one_out_reg[15]  ( .G(1'b1), .D(N975), .Q(Data_one_out[15]) );
  DLH_X1 \Data_one_out_reg[11]  ( .G(1'b1), .D(N971), .Q(Data_one_out[11]) );
  DLH_X1 \Data_one_out_reg[10]  ( .G(1'b1), .D(N970), .Q(Data_one_out[10]) );
  DLH_X1 \Data_one_out_reg[8]  ( .G(1'b1), .D(N968), .Q(Data_one_out[8]) );
  DLH_X1 \Data_one_out_reg[7]  ( .G(1'b1), .D(N967), .Q(Data_one_out[7]) );
  DLH_X1 \Data_one_out_reg[6]  ( .G(1'b1), .D(N966), .Q(Data_one_out[6]) );
  DLH_X1 \Data_one_out_reg[1]  ( .G(1'b1), .D(N961), .Q(Data_one_out[1]) );
  DLH_X1 \Data_two_out_reg[31]  ( .G(1'b1), .D(N1024), .Q(Data_two_out[31]) );
  DLH_X1 \Data_two_out_reg[30]  ( .G(1'b1), .D(N1023), .Q(Data_two_out[30]) );
  DLH_X1 \Data_two_out_reg[29]  ( .G(1'b1), .D(N1022), .Q(Data_two_out[29]) );
  DLH_X1 \Data_two_out_reg[28]  ( .G(1'b1), .D(N1021), .Q(Data_two_out[28]) );
  DLH_X1 \Data_two_out_reg[27]  ( .G(1'b1), .D(N1020), .Q(Data_two_out[27]) );
  DLH_X1 \Data_two_out_reg[26]  ( .G(1'b1), .D(N1019), .Q(Data_two_out[26]) );
  DLH_X1 \Data_two_out_reg[25]  ( .G(1'b1), .D(N1018), .Q(Data_two_out[25]) );
  DLH_X1 \Data_two_out_reg[24]  ( .G(1'b1), .D(N1017), .Q(Data_two_out[24]) );
  DLH_X1 \Data_two_out_reg[23]  ( .G(1'b1), .D(N1016), .Q(Data_two_out[23]) );
  DLH_X1 \Data_two_out_reg[22]  ( .G(1'b1), .D(N1015), .Q(Data_two_out[22]) );
  DLH_X1 \Data_two_out_reg[21]  ( .G(1'b1), .D(N1014), .Q(Data_two_out[21]) );
  DLH_X1 \Data_two_out_reg[20]  ( .G(1'b1), .D(N1013), .Q(Data_two_out[20]) );
  DLH_X1 \Data_two_out_reg[19]  ( .G(1'b1), .D(N1012), .Q(Data_two_out[19]) );
  DLH_X1 \Data_two_out_reg[18]  ( .G(1'b1), .D(N1011), .Q(Data_two_out[18]) );
  DLH_X1 \Data_two_out_reg[17]  ( .G(1'b1), .D(N1010), .Q(Data_two_out[17]) );
  DLH_X1 \Data_two_out_reg[16]  ( .G(1'b1), .D(N1009), .Q(Data_two_out[16]) );
  DLH_X1 \Data_two_out_reg[15]  ( .G(1'b1), .D(N1008), .Q(Data_two_out[15]) );
  DLH_X1 \Data_two_out_reg[14]  ( .G(1'b1), .D(N1007), .Q(Data_two_out[14]) );
  DLH_X1 \Data_two_out_reg[13]  ( .G(1'b1), .D(N1006), .Q(Data_two_out[13]) );
  DLH_X1 \Data_two_out_reg[12]  ( .G(1'b1), .D(N1005), .Q(Data_two_out[12]) );
  DLH_X1 \Data_two_out_reg[11]  ( .G(1'b1), .D(N1004), .Q(Data_two_out[11]) );
  DLH_X1 \Data_two_out_reg[10]  ( .G(1'b1), .D(N1003), .Q(Data_two_out[10]) );
  DLH_X1 \Data_two_out_reg[9]  ( .G(1'b1), .D(N1002), .Q(Data_two_out[9]) );
  DLH_X1 \Data_two_out_reg[8]  ( .G(1'b1), .D(N1001), .Q(Data_two_out[8]) );
  DLH_X1 \Data_two_out_reg[7]  ( .G(1'b1), .D(N1000), .Q(Data_two_out[7]) );
  DLH_X1 \Data_two_out_reg[6]  ( .G(1'b1), .D(N999), .Q(Data_two_out[6]) );
  DLH_X1 \Data_two_out_reg[5]  ( .G(1'b1), .D(N998), .Q(Data_two_out[5]) );
  DLH_X1 \Data_two_out_reg[4]  ( .G(1'b1), .D(N997), .Q(Data_two_out[4]) );
  DLH_X1 \Data_two_out_reg[3]  ( .G(1'b1), .D(N996), .Q(Data_two_out[3]) );
  DLH_X1 \Data_two_out_reg[2]  ( .G(1'b1), .D(N995), .Q(Data_two_out[2]) );
  DLH_X1 \Data_two_out_reg[1]  ( .G(1'b1), .D(N994), .Q(Data_two_out[1]) );
  DLH_X1 \Data_two_out_reg[0]  ( .G(1'b1), .D(N993), .Q(Data_two_out[0]) );
  DLH_X1 \Data_one_out_reg[12]  ( .G(1'b1), .D(N972), .Q(Data_one_out[12]) );
  DLH_X1 \Data_one_out_reg[0]  ( .G(1'b1), .D(N960), .Q(Data_one_out[0]) );
  DLH_X1 \Data_one_out_reg[5]  ( .G(1'b1), .D(N965), .Q(Data_one_out[5]) );
  DLH_X1 \Data_one_out_reg[17]  ( .G(1'b1), .D(N977), .Q(Data_one_out[17]) );
  DLH_X1 \Data_one_out_reg[22]  ( .G(1'b1), .D(N982), .Q(Data_one_out[22]) );
  DLH_X1 \Data_one_out_reg[24]  ( .G(1'b1), .D(N984), .Q(Data_one_out[24]) );
  DLH_X1 \Data_one_out_reg[3]  ( .G(1'b1), .D(N963), .Q(Data_one_out[3]) );
  DLH_X1 \Data_one_out_reg[2]  ( .G(1'b1), .D(N962), .Q(Data_one_out[2]) );
  DLH_X1 \Data_one_out_reg[4]  ( .G(1'b1), .D(N964), .Q(Data_one_out[4]) );
  DLH_X1 \Data_one_out_reg[9]  ( .G(1'b1), .D(N969), .Q(Data_one_out[9]) );
  DLH_X1 \Data_one_out_reg[19]  ( .G(1'b1), .D(N979), .Q(Data_one_out[19]) );
  DLH_X1 \Data_one_out_reg[18]  ( .G(1'b1), .D(N978), .Q(Data_one_out[18]) );
  DLH_X1 \Data_one_out_reg[14]  ( .G(1'b1), .D(N974), .Q(Data_one_out[14]) );
  DLH_X1 \Data_one_out_reg[13]  ( .G(1'b1), .D(N973), .Q(Data_one_out[13]) );
  DLH_X1 \Data_one_out_reg[16]  ( .G(1'b1), .D(N976), .Q(Data_one_out[16]) );
  OAI33_X1 U3389 ( .A1(n1440), .A2(n1441), .A3(n1449), .B1(n1453), .B2(n1454), 
        .B3(n1463), .ZN(n1439) );
  OAI33_X1 U3390 ( .A1(n1703), .A2(n1704), .A3(n1712), .B1(n1715), .B2(n1716), 
        .B3(n1718), .ZN(n1702) );
  OAI33_X1 U3391 ( .A1(n1776), .A2(n1777), .A3(n1779), .B1(n1780), .B2(n1781), 
        .B3(n1782), .ZN(n1774) );
  NAND3_X1 U3392 ( .A1(n1828), .A2(n1830), .A3(n1831), .ZN(N988) );
  OAI33_X1 U3393 ( .A1(n1843), .A2(n1844), .A3(n1845), .B1(n1848), .B2(n1849), 
        .B3(n1850), .ZN(n1842) );
  NAND3_X1 U3394 ( .A1(n2095), .A2(n2096), .A3(n2097), .ZN(N984) );
  OAI33_X1 U3395 ( .A1(n2104), .A2(n2105), .A3(n2106), .B1(n2107), .B2(n2108), 
        .B3(n2109), .ZN(n2101) );
  NAND3_X1 U3396 ( .A1(n2158), .A2(n2159), .A3(n2160), .ZN(N982) );
  OAI33_X1 U3397 ( .A1(n2165), .A2(n2166), .A3(n2167), .B1(n2168), .B2(n2169), 
        .B3(n2170), .ZN(n2164) );
  NAND3_X1 U3398 ( .A1(n2234), .A2(n2235), .A3(n2236), .ZN(N978) );
  OAI33_X1 U3399 ( .A1(n2241), .A2(n2242), .A3(n2243), .B1(n2244), .B2(n2245), 
        .B3(n2246), .ZN(n2240) );
  NAND3_X1 U3400 ( .A1(n2252), .A2(n2253), .A3(n2254), .ZN(N977) );
  OAI33_X1 U3401 ( .A1(n2258), .A2(n2259), .A3(n2260), .B1(n2261), .B2(n2262), 
        .B3(n2263), .ZN(n2257) );
  NAND3_X1 U3402 ( .A1(n2305), .A2(n2306), .A3(n2307), .ZN(N974) );
  OAI33_X1 U3403 ( .A1(n2312), .A2(n2313), .A3(n2314), .B1(n2315), .B2(n2316), 
        .B3(n2317), .ZN(n2311) );
  NAND3_X1 U3404 ( .A1(n2323), .A2(n2324), .A3(n2325), .ZN(N973) );
  NAND3_X1 U3405 ( .A1(n2434), .A2(n14844), .A3(n2435), .ZN(n2433) );
  NAND3_X1 U3406 ( .A1(n2452), .A2(n2453), .A3(n2454), .ZN(N966) );
  NAND3_X1 U3407 ( .A1(n2469), .A2(n2470), .A3(n2471), .ZN(N965) );
  OAI33_X1 U3408 ( .A1(n2476), .A2(n2477), .A3(n2478), .B1(n2479), .B2(n2480), 
        .B3(n2481), .ZN(n2475) );
  NAND3_X1 U3409 ( .A1(n2487), .A2(n2488), .A3(n2489), .ZN(N964) );
  NAND3_X1 U3410 ( .A1(n14844), .A2(n14619), .A3(n2543), .ZN(n2542) );
  NAND3_X1 U3411 ( .A1(n2560), .A2(n2561), .A3(n2562), .ZN(N960) );
  OAI33_X1 U3412 ( .A1(n2568), .A2(n2569), .A3(n2570), .B1(n2571), .B2(n2572), 
        .B3(n2573), .ZN(n2567) );
  NAND3_X1 U3413 ( .A1(Read_one_address[2]), .A2(n15303), .A3(
        Read_one_address[4]), .ZN(n1471) );
  NAND3_X1 U3414 ( .A1(Read_one_address[3]), .A2(Read_one_address[2]), .A3(
        Read_one_address[4]), .ZN(n1656) );
  NAND3_X1 U3415 ( .A1(Read_one_address[2]), .A2(n15347), .A3(
        Read_one_address[3]), .ZN(n1639) );
  NAND3_X1 U3416 ( .A1(Read_one_address[3]), .A2(n15301), .A3(
        Read_one_address[4]), .ZN(n1662) );
  XOR2_X1 U3417 ( .A(Write_address[3]), .B(Read_one_address[3]), .Z(n2585) );
  XOR2_X1 U3418 ( .A(Write_address[0]), .B(n15278), .Z(n2584) );
  XOR2_X1 U3419 ( .A(Write_address[4]), .B(Read_one_address[4]), .Z(n2583) );
  XOR2_X1 U3420 ( .A(n15311), .B(Read_one_address[1]), .Z(n2581) );
  XOR2_X1 U3421 ( .A(n15301), .B(Write_address[2]), .Z(n2579) );
  XOR2_X1 U3422 ( .A(Write_address[3]), .B(Read_two_address[3]), .Z(n3054) );
  XOR2_X1 U3423 ( .A(Write_address[0]), .B(Read_two_address[0]), .Z(n3052) );
  XOR2_X1 U3424 ( .A(Write_address[4]), .B(Read_two_address[4]), .Z(n3051) );
  XOR2_X1 U3425 ( .A(n15282), .B(Write_address[2]), .Z(n3049) );
  XOR2_X1 U3426 ( .A(n15281), .B(Write_address[1]), .Z(n3048) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n2073), .CK(CK), .RN(n14606), .Q(n15485), .QN(n9444) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3760), .CK(CK), .RN(n14605), .Q(n15479), .QN(n3383) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n2066), .CK(CK), .RN(n14607), .Q(n15488), .QN(n9445) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n2063), .CK(CK), .RN(n14606), .Q(n15492), .QN(n9443) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3762), .CK(CK), .RN(n14605), .Q(n15481), 
        .QN(n3594) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n2015), .CK(CK), .RN(n14607), .Q(n15354), .QN(n9591) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n2014), .CK(CK), .RN(n14606), .Q(n15355), .QN(n9590) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n2010), .CK(CK), .RN(n14605), .Q(n15356), .QN(n9586) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n2008), .CK(CK), .RN(n14607), .Q(n15357), .QN(n9587) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n2004), .CK(CK), .RN(n14606), .Q(n15358), .QN(n9585) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n1991), .CK(CK), .RN(n14605), .Q(n15359), 
        .QN(n9588) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n1986), .CK(CK), .RN(n14607), .Q(n15361), 
        .QN(n9589) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n1833), .CK(CK), .RN(n14606), .Q(n15374), 
        .QN(n7813) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n1751), .CK(CK), .RN(n14605), .Q(n15376), .QN(n9580) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n1742), .CK(CK), .RN(n14607), .Q(n15377), .QN(n9581) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n1741), .CK(CK), .RN(n14606), .Q(n15378), .QN(n9579) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n1738), .CK(CK), .RN(n14605), .Q(n15462), 
        .QN(n9576) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n1733), .CK(CK), .RN(n14607), .Q(n15464), 
        .QN(n9577) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n1591), .CK(CK), .RN(n14606), .Q(n15465), .QN(n9469) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n1582), .CK(CK), .RN(n14605), .Q(n15466), .QN(n9468) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n1581), .CK(CK), .RN(n14607), .Q(n15467), .QN(n9467) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n1203), .CK(CK), .RN(n14606), .Q(n15398), 
        .QN(n9433) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n1200), .CK(CK), .RN(n14605), .Q(n15450), 
        .QN(n9583) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n1193), .CK(CK), .RN(n14607), .Q(n15478), 
        .QN(n9566) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n1185), .CK(CK), .RN(n14606), .Q(n15460), 
        .QN(n8080) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n1184), .CK(CK), .RN(n14605), .Q(n15461), 
        .QN(n8079) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3483), .CK(CK), .RN(n14607), .Q(n15407), 
        .QN(n3362) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3492), .CK(CK), .RN(n14606), .Q(n15410), 
        .QN(n3356) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3587), .CK(CK), .RN(n14605), .Q(n15411), 
        .QN(n3240) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3484), .CK(CK), .RN(n14607), .Q(n15412), 
        .QN(n3337) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n1175), .CK(CK), .RN(n14606), .Q(n15413), 
        .QN(n8100) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3485), .CK(CK), .RN(n14605), .Q(n15414), 
        .QN(n3358) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3486), .CK(CK), .RN(n14607), .Q(n15415), 
        .QN(n3333) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3588), .CK(CK), .RN(n14606), .Q(n15416), 
        .QN(n3329) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n1166), .CK(CK), .RN(n14605), .Q(n15417), 
        .QN(n7831) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n1165), .CK(CK), .RN(n14607), .Q(n15418), 
        .QN(n7830) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3488), .CK(CK), .RN(n14606), .Q(n15421), 
        .QN(n3335) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3489), .CK(CK), .RN(n14605), .Q(n15422), 
        .QN(n3381) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3490), .CK(CK), .RN(n14607), .Q(n15423), 
        .QN(n3354) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3491), .CK(CK), .RN(n14606), .Q(n15425), 
        .QN(n3360) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n3735), .CK(CK), .RN(n14605), .QN(n3681)
         );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n3736), .CK(CK), .RN(n14607), .QN(n3680)
         );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n3737), .CK(CK), .RN(n14606), .QN(n3682)
         );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n3781), .CK(CK), .RN(n14605), .QN(n3379)
         );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n3782), .CK(CK), .RN(n14607), .QN(n3375)
         );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n3783), .CK(CK), .RN(n14606), .QN(n3374)
         );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n3784), .CK(CK), .RN(n14605), .QN(n3373)
         );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n3785), .CK(CK), .RN(n14607), .QN(n3372)
         );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n1815), .CK(CK), .RN(n14606), .QN(n9723) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n1806), .CK(CK), .RN(n14605), .QN(n9722) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n1805), .CK(CK), .RN(n14607), .QN(n9721) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n1936), .CK(CK), .RN(n14606), .Q(n15463), .QN(n9450) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n1527), .CK(CK), .RN(n14605), .Q(n15380), .QN(n9575) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n1518), .CK(CK), .RN(n14607), .Q(n15381), .QN(n9573) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n1517), .CK(CK), .RN(n14606), .Q(n15382), .QN(n9574) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n1407), .CK(CK), .RN(n14605), .Q(n15446), 
        .QN(n9438) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n3778), .CK(CK), .RN(n14607), .Q(n15447), 
        .QN(n3382) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n1386), .CK(CK), .RN(n14606), .Q(n15448), 
        .QN(n9503) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n1385), .CK(CK), .RN(n14605), .Q(n15449), 
        .QN(n9502) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n2064), .CK(CK), .RN(n14607), .Q(n15480), .QN(n9341) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n1217), .CK(CK), .RN(n14606), .Q(n15453), 
        .QN(n9435) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n1216), .CK(CK), .RN(n14605), .Q(n15454), 
        .QN(n9434) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3754), .CK(CK), .RN(n14607), .Q(n15403), 
        .QN(n3365) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3786), .CK(CK), .RN(n14606), .Q(n15379), 
        .QN(n3640) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n2043), .CK(CK), .RN(n14605), .QN(n9739) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n2037), .CK(CK), .RN(n14607), .QN(n9735) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n2033), .CK(CK), .RN(n14606), .QN(n9734) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3739), .CK(CK), .RN(n14605), .QN(n3348)
         );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3743), .CK(CK), .RN(n14607), .QN(n3347)
         );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3744), .CK(CK), .RN(n14606), .QN(n3346)
         );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n1987), .CK(CK), .RN(n14605), .Q(n15360), 
        .QN(n9592) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3532), .CK(CK), .RN(n14607), .Q(n15457), .QN(n3224) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3533), .CK(CK), .RN(n14606), .Q(n15458), .QN(n3229) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3535), .CK(CK), .RN(n14605), .Q(n15368), .QN(n3228) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3536), .CK(CK), .RN(n14607), .Q(n15369), .QN(n3227) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3537), .CK(CK), .RN(n14606), .Q(n15370), .QN(n3226) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3541), .CK(CK), .RN(n14605), .Q(n15371), .QN(n3225) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3545), .CK(CK), .RN(n14607), .Q(n15372), .QN(n3203) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3548), .CK(CK), .RN(n14606), .Q(n15373), .QN(n3310) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3553), .CK(CK), .RN(n14605), .Q(n15375), 
        .QN(n3311) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3748), .CK(CK), .RN(n14607), .Q(n15393), 
        .QN(n3371) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3749), .CK(CK), .RN(n14606), .Q(n15394), 
        .QN(n3370) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3750), .CK(CK), .RN(n14605), .Q(n15395), 
        .QN(n3369) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3751), .CK(CK), .RN(n14607), .Q(n15397), 
        .QN(n3368) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3752), .CK(CK), .RN(n14606), .Q(n15399), 
        .QN(n3367) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3753), .CK(CK), .RN(n14605), .Q(n15402), 
        .QN(n3366) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n1192), .CK(CK), .RN(n14607), .Q(n15404), 
        .QN(n9449) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n1190), .CK(CK), .RN(n14606), .Q(n15405), 
        .QN(n9448) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3755), .CK(CK), .RN(n14605), .Q(n15451), 
        .QN(n3364) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3756), .CK(CK), .RN(n14607), .Q(n15406), 
        .QN(n3363) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n1181), .CK(CK), .RN(n14606), .Q(n15408), 
        .QN(n8086) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n1180), .CK(CK), .RN(n14605), .Q(n15409), 
        .QN(n8085) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n1164), .CK(CK), .RN(n14607), .Q(n15419), 
        .QN(n7822) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n1156), .CK(CK), .RN(n14606), .Q(n15424), 
        .QN(n7821) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n3934), .CK(CK), .RN(n14605), .Q(n15482), 
        .QN(n3929) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3590), .CK(CK), .RN(n14607), .Q(n15452), 
        .QN(n3242) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n3765), .CK(CK), .RN(n14606), .Q(n15362), .QN(n3654) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n3766), .CK(CK), .RN(n14605), .Q(n15363), .QN(n3656) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n3767), .CK(CK), .RN(n14607), .Q(n15364), .QN(n3653) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n3769), .CK(CK), .RN(n14606), .Q(n15365), .QN(n3657) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n3772), .CK(CK), .RN(n14605), .Q(n15366), 
        .QN(n3658) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n3773), .CK(CK), .RN(n14607), .Q(n15367), 
        .QN(n3655) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3779), .CK(CK), .RN(n14606), .Q(n15468), 
        .QN(n3724) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3780), .CK(CK), .RN(n14605), .Q(n15469), 
        .QN(n3725) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3757), .CK(CK), .RN(n14607), .Q(n15483), .QN(n3642) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3758), .CK(CK), .RN(n14606), .Q(n15484), .QN(n3643) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3759), .CK(CK), .RN(n14605), .Q(n15486), .QN(n3361) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3935), .CK(CK), .RN(n14607), .Q(n15491), .QN(n3932) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3761), .CK(CK), .RN(n14606), .Q(n15487), .QN(n3359) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3936), .CK(CK), .RN(n14605), .Q(n15493), .QN(n3931) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3937), .CK(CK), .RN(n14607), .Q(n15494), .QN(n3930) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3763), .CK(CK), .RN(n14606), .Q(n15489), 
        .QN(n3357) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3764), .CK(CK), .RN(n14605), .Q(n15490), 
        .QN(n3355) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n2049), .CK(CK), .RN(n14607), .Q(n15348), .QN(n9738) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n2048), .CK(CK), .RN(n14606), .Q(n15349), .QN(n9737) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n2045), .CK(CK), .RN(n14605), .Q(n15350), .QN(n9740) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n2044), .CK(CK), .RN(n14607), .Q(n15351), .QN(n9736) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n2028), .CK(CK), .RN(n14606), .Q(n15352), .QN(n9732) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n2020), .CK(CK), .RN(n14605), .Q(n15353), 
        .QN(n9733) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3549), .CK(CK), .RN(n14607), .Q(n15459), 
        .QN(n3208) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n1482), .CK(CK), .RN(n14606), .Q(n15445), 
        .QN(n9725) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n1470), .CK(CK), .RN(n14605), .Q(n15383), .QN(n9451) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n1466), .CK(CK), .RN(n14607), .Q(n15384), .QN(n9594) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n1464), .CK(CK), .RN(n14606), .Q(n15385), .QN(n9595) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3731), .CK(CK), .RN(n14605), .Q(n15386), .QN(n3631) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n1462), .CK(CK), .RN(n14607), .Q(n15387), .QN(n9439) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n1460), .CK(CK), .RN(n14606), .Q(n15388), .QN(n9593) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3732), .CK(CK), .RN(n14605), .Q(n15389), .QN(n3630) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3733), .CK(CK), .RN(n14607), .Q(n15390), .QN(n3629) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n1447), .CK(CK), .RN(n14606), .Q(n15391), 
        .QN(n9596) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n1442), .CK(CK), .RN(n14605), .Q(n15392), 
        .QN(n9597) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n1555), .CK(CK), .RN(n14607), .QN(n9571) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n1544), .CK(CK), .RN(n14606), .QN(n9572)
         );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n1542), .CK(CK), .RN(n14605), .QN(n9570)
         );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3591), .CK(CK), .RN(n14607), .Q(n15420), 
        .QN(n3147) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n2007), .CK(CK), .RN(n14606), .Q(n15470), .QN(n9441) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n2006), .CK(CK), .RN(n14605), .Q(n15471), .QN(n9891) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n1998), .CK(CK), .RN(n14607), .Q(n15472), .QN(n9442) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n1997), .CK(CK), .RN(n14606), .Q(n15473), .QN(n9440) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n3768), .CK(CK), .RN(n14605), .Q(n15474), .QN(n3353) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n1974), .CK(CK), .RN(n14607), .Q(n15475), .QN(n9506) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n3770), .CK(CK), .RN(n14606), .Q(n15476), .QN(n3352) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n3771), .CK(CK), .RN(n14605), .Q(n15477), .QN(n3351) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n1207), .CK(CK), .RN(n14607), .Q(n15396), 
        .QN(n9446) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n1198), .CK(CK), .RN(n14606), .Q(n15400), 
        .QN(n9582) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n1197), .CK(CK), .RN(n14605), .Q(n15401), 
        .QN(n9447) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n3980), .CK(CK), .RN(n14607), .Q(n15499), 
        .QN(n3979) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n15305), .CK(CK), .RN(n14606), .Q(n3245) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n15306), .CK(CK), .RN(n14605), .Q(n3258) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n15307), .CK(CK), .RN(n14607), .Q(n3244) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n15308), .CK(CK), .RN(n14606), .Q(n3243) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n15309), .CK(CK), .RN(n14605), .Q(n3239)
         );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n15310), .CK(CK), .RN(n14607), .Q(n3236)
         );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n3600), .CK(CK), .RN(n14606), .QN(n16141) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n3601), .CK(CK), .RN(n14605), .QN(n16142) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n3602), .CK(CK), .RN(n14607), .QN(n16143) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n3603), .CK(CK), .RN(n14606), .QN(n16144) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n1267), .CK(CK), .RN(n14605), .QN(n16145) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n1264), .CK(CK), .RN(n14607), .QN(n16068) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n1259), .CK(CK), .RN(n14606), .QN(n16069)
         );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n1256), .CK(CK), .RN(n14605), .QN(n16070)
         );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n3604), .CK(CK), .RN(n14607), .QN(n16146)
         );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n1254), .CK(CK), .RN(n14606), .QN(n16071)
         );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n3605), .CK(CK), .RN(n14605), .QN(n16147)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n1939), .CK(CK), .RN(n14607), .QN(
        n15735) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n1928), .CK(CK), .RN(n14606), .QN(n15736) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n1926), .CK(CK), .RN(n14605), .QN(n15737) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n1615), .CK(CK), .RN(n14607), .QN(
        n15746) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n1406), .CK(CK), .RN(n14606), .QN(n15608) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n1402), .CK(CK), .RN(n14605), .QN(n15609) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n1400), .CK(CK), .RN(n14607), .QN(n15610) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n1396), .CK(CK), .RN(n14606), .QN(n15611) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n1383), .CK(CK), .RN(n14605), .QN(n15612)
         );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n1378), .CK(CK), .RN(n14607), .QN(n15614)
         );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n3563), .CK(CK), .RN(n14606), .QN(n15933) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n3564), .CK(CK), .RN(n14605), .QN(n15934) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n3568), .CK(CK), .RN(n14607), .QN(n16078) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n3569), .CK(CK), .RN(n14606), .QN(n16079) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n3570), .CK(CK), .RN(n14605), .QN(n16080) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n1253), .CK(CK), .RN(n14607), .QN(n16082)
         );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n1807), .CK(CK), .RN(n14606), .QN(
        n15729) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n1609), .CK(CK), .RN(n14605), .QN(n15543) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n1931), .CK(CK), .RN(n14607), .QN(n15563) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3528), .CK(CK), .RN(n14606), .QN(n16043) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3529), .CK(CK), .RN(n14605), .QN(n16044) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n1822), .CK(CK), .RN(n14607), .QN(
        n15588) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n1821), .CK(CK), .RN(n14606), .QN(
        n15620) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n1820), .CK(CK), .RN(n14605), .QN(
        n15621) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n1818), .CK(CK), .RN(n14607), .QN(
        n15589) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n1816), .CK(CK), .RN(n14606), .QN(
        n15590) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n1812), .CK(CK), .RN(n14605), .QN(
        n15591) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n1804), .CK(CK), .RN(n14607), .QN(
        n15622) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n1799), .CK(CK), .RN(n14606), .QN(n15594) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n1796), .CK(CK), .RN(n14605), .QN(n15623) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n1794), .CK(CK), .RN(n14607), .QN(n15596) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n1531), .CK(CK), .RN(n14606), .QN(
        n15762) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n1525), .CK(CK), .RN(n14605), .QN(
        n15763) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n1521), .CK(CK), .RN(n14607), .QN(
        n15764) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n1509), .CK(CK), .RN(n14606), .QN(n15767) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n1405), .CK(CK), .RN(n14605), .QN(n15441) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n1404), .CK(CK), .RN(n14607), .QN(n15442) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n1388), .CK(CK), .RN(n14606), .QN(n15443) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n1381), .CK(CK), .RN(n14605), .QN(n15685)
         );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n1380), .CK(CK), .RN(n14607), .QN(n15444)
         );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n1913), .CK(CK), .RN(n14606), .QN(
        n16061) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n1906), .CK(CK), .RN(n14605), .QN(
        n16064) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n1891), .CK(CK), .RN(n14607), .QN(n15921) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n1785), .CK(CK), .RN(n14606), .QN(
        n16024) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n1778), .CK(CK), .RN(n14605), .QN(
        n16026) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n1263), .CK(CK), .RN(n14607), .QN(n15922) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n1251), .CK(CK), .RN(n14606), .QN(n16140)
         );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n1921), .CK(CK), .RN(n14605), .QN(
        n15923) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n1920), .CK(CK), .RN(n14607), .QN(
        n15924) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n1915), .CK(CK), .RN(n14606), .QN(
        n16018) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n1909), .CK(CK), .RN(n14605), .QN(
        n16019) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n1905), .CK(CK), .RN(n14607), .QN(
        n16020) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n1893), .CK(CK), .RN(n14606), .QN(n16022) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n1391), .CK(CK), .RN(n14605), .QN(n15633) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n1379), .CK(CK), .RN(n14607), .QN(n15613)
         );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n1546), .CK(CK), .RN(n14606), .QN(n15669) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n1545), .CK(CK), .RN(n14605), .QN(n15670) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n1795), .CK(CK), .RN(n14607), .QN(n15730) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3774), .CK(CK), .RN(n14606), .QN(
        n15552) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3776), .CK(CK), .RN(n14605), .QN(
        n15555) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3512), .CK(CK), .RN(n14607), .QN(
        n16012) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3513), .CK(CK), .RN(n14606), .QN(
        n16013) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n1533), .CK(CK), .RN(n14605), .QN(
        n15776) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n1532), .CK(CK), .RN(n14607), .QN(
        n15777) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n1516), .CK(CK), .RN(n14606), .QN(
        n15778) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n1508), .CK(CK), .RN(n14605), .QN(n15779) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n1925), .CK(CK), .RN(n14607), .QN(n15508) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n1923), .CK(CK), .RN(n14606), .QN(n15532) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3527), .CK(CK), .RN(n14605), .QN(n16089) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n1803), .CK(CK), .RN(n14607), .QN(n15671) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n2046), .CK(CK), .RN(n14606), .QN(
        n15893) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n2042), .CK(CK), .RN(n14605), .QN(
        n15894) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n2040), .CK(CK), .RN(n14607), .QN(
        n15895) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n2036), .CK(CK), .RN(n14606), .QN(
        n15896) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n2035), .CK(CK), .RN(n14605), .QN(
        n15897) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n2032), .CK(CK), .RN(n14607), .QN(
        n15898) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n2027), .CK(CK), .RN(n14606), .QN(n15900) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n2024), .CK(CK), .RN(n14605), .QN(n15901) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n2023), .CK(CK), .RN(n14607), .QN(n15902) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n2022), .CK(CK), .RN(n14606), .QN(n15903) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n2018), .CK(CK), .RN(n14605), .QN(n15904) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n3395), .CK(CK), .RN(n14607), .QN(
        n15927) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n3396), .CK(CK), .RN(n14606), .QN(
        n15928) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n3397), .CK(CK), .RN(n14605), .QN(
        n16120) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n3581), .CK(CK), .RN(n14607), .QN(
        n16121) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n3404), .CK(CK), .RN(n14606), .QN(
        n16122) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n3408), .CK(CK), .RN(n14605), .QN(
        n15929) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n3415), .CK(CK), .RN(n14607), .QN(n16123) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n3416), .CK(CK), .RN(n14606), .QN(n15930) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n1675), .CK(CK), .RN(n14605), .QN(n16038) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n1674), .CK(CK), .RN(n14607), .QN(n15953) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n1673), .CK(CK), .RN(n14606), .QN(n15954) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n1669), .CK(CK), .RN(n14605), .QN(n16095) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3738), .CK(CK), .RN(n14607), .QN(n15908) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3740), .CK(CK), .RN(n14606), .QN(n15910) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3734), .CK(CK), .RN(n14605), .QN(n15863) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n1695), .CK(CK), .RN(n14607), .QN(
        n16124) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n1687), .CK(CK), .RN(n14606), .QN(
        n16125) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n1678), .CK(CK), .RN(n14605), .QN(
        n16126) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n1677), .CK(CK), .RN(n14607), .QN(
        n16127) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n1551), .CK(CK), .RN(n14606), .QN(
        n15581) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n1473), .CK(CK), .RN(n14605), .QN(
        n15843) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n1472), .CK(CK), .RN(n14607), .QN(
        n15844) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n1469), .CK(CK), .RN(n14606), .QN(
        n15659) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n1468), .CK(CK), .RN(n14605), .QN(
        n15660) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n1467), .CK(CK), .RN(n14607), .QN(
        n15661) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n1461), .CK(CK), .RN(n14606), .QN(
        n15662) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n1457), .CK(CK), .RN(n14605), .QN(
        n15663) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n1452), .CK(CK), .RN(n14607), .QN(
        n15664) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n1445), .CK(CK), .RN(n14606), .QN(n15665) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n1444), .CK(CK), .RN(n14605), .QN(n15666) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n1443), .CK(CK), .RN(n14607), .QN(n15667) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n1245), .CK(CK), .RN(n14606), .QN(n15823) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n1244), .CK(CK), .RN(n14605), .QN(n15824) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n1243), .CK(CK), .RN(n14607), .QN(n15825) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n1237), .CK(CK), .RN(n14606), .QN(n15826) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n1233), .CK(CK), .RN(n14605), .QN(n15827) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n1228), .CK(CK), .RN(n14607), .QN(n15828) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3745), .CK(CK), .RN(n14606), .QN(n15769)
         );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n1226), .CK(CK), .RN(n14605), .QN(n15829)
         );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3746), .CK(CK), .RN(n14607), .QN(n15770)
         );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3747), .CK(CK), .RN(n14606), .QN(n15771)
         );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n1221), .CK(CK), .RN(n14605), .QN(n15831)
         );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n1220), .CK(CK), .RN(n14607), .QN(n15832)
         );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n1219), .CK(CK), .RN(n14606), .QN(n15852)
         );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n2041), .CK(CK), .RN(n14605), .QN(
        n15917) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n2034), .CK(CK), .RN(n14607), .QN(
        n15918) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n2019), .CK(CK), .RN(n14606), .QN(n15912) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n1238), .CK(CK), .RN(n14605), .QN(n15905) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n1455), .CK(CK), .RN(n14607), .QN(
        n15694) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3425), .CK(CK), .RN(n14606), .QN(
        n16296) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n1693), .CK(CK), .RN(n14605), .QN(
        n15974) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n1692), .CK(CK), .RN(n14607), .QN(
        n15975) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n1686), .CK(CK), .RN(n14606), .QN(
        n15961) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n1676), .CK(CK), .RN(n14605), .QN(
        n15977) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n1668), .CK(CK), .RN(n14607), .QN(n15980) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n1567), .CK(CK), .RN(n14606), .QN(
        n15510) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n1448), .CK(CK), .RN(n14605), .QN(n15695) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n1446), .CK(CK), .RN(n14607), .QN(n15696) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n1246), .CK(CK), .RN(n14606), .QN(n15886) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n1242), .CK(CK), .RN(n14605), .QN(n15887) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n1240), .CK(CK), .RN(n14607), .QN(n15888) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n1236), .CK(CK), .RN(n14606), .QN(n15889) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n1223), .CK(CK), .RN(n14605), .QN(n15890)
         );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n1218), .CK(CK), .RN(n14607), .QN(n15891)
         );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n1721), .CK(CK), .RN(n14606), .QN(
        n16264) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n1714), .CK(CK), .RN(n14605), .QN(
        n16265) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3742), .CK(CK), .RN(n14607), .QN(n15851) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n2021), .CK(CK), .RN(n14606), .QN(n15789) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n1705), .CK(CK), .RN(n14605), .QN(n16244) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n1689), .CK(CK), .RN(n14607), .QN(
        n16014) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n1682), .CK(CK), .RN(n14606), .QN(
        n16015) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n1679), .CK(CK), .RN(n14605), .QN(
        n16037) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n1566), .CK(CK), .RN(n14607), .QN(
        n15522) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n1562), .CK(CK), .RN(n14606), .QN(
        n15524) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n1560), .CK(CK), .RN(n14605), .QN(
        n15525) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n1556), .CK(CK), .RN(n14607), .QN(
        n15527) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n1543), .CK(CK), .RN(n14606), .QN(n15529) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n1538), .CK(CK), .RN(n14605), .QN(n15530) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n1450), .CK(CK), .RN(n14607), .QN(n15701) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n1949), .CK(CK), .RN(n14606), .Q(n9340), 
        .QN(n15634) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n1948), .CK(CK), .RN(n14605), .Q(n9339), 
        .QN(n15635) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n1947), .CK(CK), .RN(n14607), .Q(n3316), 
        .QN(n15615) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n1941), .CK(CK), .RN(n14606), .Q(n3314), 
        .QN(n15616) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n1937), .CK(CK), .RN(n14605), .Q(n3308), 
        .QN(n15617) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3777), .CK(CK), .RN(n14607), .Q(n3917), 
        .QN(n15587) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n1932), .CK(CK), .RN(n14606), .Q(n9338), 
        .QN(n15636) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n1930), .CK(CK), .RN(n14605), .Q(n3301), 
        .QN(n15618) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n1929), .CK(CK), .RN(n14607), .Q(n3300), 
        .QN(n15619) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n1924), .CK(CK), .RN(n14606), .Q(n9337), 
        .QN(n15637) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3517), .CK(CK), .RN(n14605), .Q(n3698), 
        .QN(n16035) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3520), .CK(CK), .RN(n14607), .Q(n3699), 
        .QN(n16036) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3523), .CK(CK), .RN(n14606), .Q(n3697), 
        .QN(n16041) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n1797), .CK(CK), .RN(n14605), .Q(n3378), 
        .QN(n15535) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n3410), .CK(CK), .RN(n14607), .Q(n3273), 
        .QN(n15951) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n3411), .CK(CK), .RN(n14606), .Q(n3272), 
        .QN(n15952) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3728), .CK(CK), .RN(n14605), .Q(n3969), 
        .QN(n15430) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3729), .CK(CK), .RN(n14607), .Q(n3968), 
        .QN(n15431) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n1817), .CK(CK), .RN(n14606), .Q(n3855), 
        .QN(n15565) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n1810), .CK(CK), .RN(n14605), .Q(n3839), 
        .QN(n15566) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n1631), .CK(CK), .RN(n14607), .Q(n3340), 
        .QN(n15559) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n1629), .CK(CK), .RN(n14606), .Q(n3667), 
        .QN(n15639) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n1628), .CK(CK), .RN(n14605), .Q(n3138), 
        .QN(n15640) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n1627), .CK(CK), .RN(n14607), .Q(n3669), 
        .QN(n15641) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n1621), .CK(CK), .RN(n14606), .Q(n3137), 
        .QN(n15642) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n1617), .CK(CK), .RN(n14605), .Q(n3136), 
        .QN(n15643) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n1616), .CK(CK), .RN(n14607), .Q(n3826), 
        .QN(n15738) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n1612), .CK(CK), .RN(n14606), .Q(n3671), 
        .QN(n15644) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n1611), .CK(CK), .RN(n14605), .Q(n3819), 
        .QN(n15739) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n1610), .CK(CK), .RN(n14607), .Q(n3866), 
        .QN(n15597) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n1605), .CK(CK), .RN(n14606), .Q(n3858), 
        .QN(n15753) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n1604), .CK(CK), .RN(n14605), .Q(n3209), 
        .QN(n15558) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n1603), .CK(CK), .RN(n14607), .Q(n3854), 
        .QN(n15747) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n3565), .CK(CK), .RN(n14606), .Q(n3299), 
        .QN(n16139) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n1271), .CK(CK), .RN(n14605), .Q(n3332), 
        .QN(n16164) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n1270), .CK(CK), .RN(n14607), .Q(n9643), 
        .QN(n16067) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n1262), .CK(CK), .RN(n14606), .Q(n3330), 
        .QN(n16165) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n1261), .CK(CK), .RN(n14605), .Q(n3328), 
        .QN(n16166) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n1886), .CK(CK), .RN(n14607), .Q(n3304), 
        .QN(n16105) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n1882), .CK(CK), .RN(n14606), .Q(n3303), 
        .QN(n16109) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n1880), .CK(CK), .RN(n14605), .Q(n3692), 
        .QN(n16110) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n1876), .CK(CK), .RN(n14607), .Q(n3693), 
        .QN(n16112) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3522), .CK(CK), .RN(n14606), .Q(n3297), 
        .QN(n16040) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n1863), .CK(CK), .RN(n14605), .Q(n3344), 
        .QN(n16116) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n1858), .CK(CK), .RN(n14607), .Q(n3341), 
        .QN(n16119) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n1802), .CK(CK), .RN(n14606), .Q(n3194), 
        .QN(n15672) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n1801), .CK(CK), .RN(n14605), .Q(n3193), 
        .QN(n15673) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3775), .CK(CK), .RN(n14607), .Q(n3961), 
        .QN(n15456) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3526), .CK(CK), .RN(n14606), .Q(n3295), 
        .QN(n16088) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n1808), .CK(CK), .RN(n14605), .Q(n3956), 
        .QN(n15560) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n1811), .CK(CK), .RN(n14607), .Q(n3928), 
        .QN(n15592) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n1800), .CK(CK), .RN(n14606), .Q(n3927), 
        .QN(n15593) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n1798), .CK(CK), .RN(n14605), .Q(n3926), 
        .QN(n15595) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n1819), .CK(CK), .RN(n14607), .Q(n3795), 
        .QN(n15726) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n1813), .CK(CK), .RN(n14606), .Q(n3702), 
        .QN(n15727) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n1809), .CK(CK), .RN(n14605), .Q(n3670), 
        .QN(n15728) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n1633), .CK(CK), .RN(n14607), .Q(n3271), 
        .QN(n15561) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n1632), .CK(CK), .RN(n14606), .Q(n3343), 
        .QN(n15562) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n1608), .CK(CK), .RN(n14605), .Q(n3864), 
        .QN(n15740) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n1606), .CK(CK), .RN(n14607), .Q(n3861), 
        .QN(n15741) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n2026), .CK(CK), .RN(n14606), .Q(n3633), 
        .QN(n15787) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n2025), .CK(CK), .RN(n14605), .Q(n3632), 
        .QN(n15788) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n1711), .CK(CK), .RN(n14607), .Q(n3093), 
        .QN(n16184) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3431), .CK(CK), .RN(n14606), .Q(n3709), 
        .QN(n16090) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3432), .CK(CK), .RN(n14605), .Q(n3159), 
        .QN(n16091) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3433), .CK(CK), .RN(n14607), .Q(n3158), 
        .QN(n16092) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3434), .CK(CK), .RN(n14606), .Q(n3156), 
        .QN(n16093) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3437), .CK(CK), .RN(n14605), .Q(n3153), 
        .QN(n16094) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3439), .CK(CK), .RN(n14607), .Q(n3711), 
        .QN(n16096) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n1569), .CK(CK), .RN(n14606), .Q(n3660), 
        .QN(n15520) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n1568), .CK(CK), .RN(n14605), .Q(n3659), 
        .QN(n15521) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n1539), .CK(CK), .RN(n14607), .Q(n3853), 
        .QN(n15579) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n1465), .CK(CK), .RN(n14606), .Q(n3833), 
        .QN(n15724) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n1458), .CK(CK), .RN(n14605), .Q(n3933), 
        .QN(n15725) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n1535), .CK(CK), .RN(n14607), .Q(n9347), 
        .QN(n15702) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n1534), .CK(CK), .RN(n14606), .Q(n9796), 
        .QN(n15703) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n1530), .CK(CK), .RN(n14605), .Q(n9795), 
        .QN(n15704) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n1528), .CK(CK), .RN(n14607), .Q(n9794), 
        .QN(n15705) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n1524), .CK(CK), .RN(n14606), .Q(n9793), 
        .QN(n15706) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n1523), .CK(CK), .RN(n14605), .Q(n9789), 
        .QN(n15707) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n1511), .CK(CK), .RN(n14607), .Q(n9792), 
        .QN(n15711) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n1507), .CK(CK), .RN(n14606), .Q(n3916), 
        .QN(n15775) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n1506), .CK(CK), .RN(n14605), .Q(n9791), 
        .QN(n15713) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n1401), .CK(CK), .RN(n14607), .Q(n3914), 
        .QN(n15495) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n1394), .CK(CK), .RN(n14606), .Q(n3886), 
        .QN(n15496) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n1565), .CK(CK), .RN(n14605), .Q(n3922), 
        .QN(n15500) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n1564), .CK(CK), .RN(n14607), .Q(n3921), 
        .QN(n15501) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n1563), .CK(CK), .RN(n14606), .Q(n3920), 
        .QN(n15523) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n1557), .CK(CK), .RN(n14605), .Q(n3891), 
        .QN(n15526) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n1553), .CK(CK), .RN(n14607), .Q(n3883), 
        .QN(n15528) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n1548), .CK(CK), .RN(n14606), .Q(n3951), 
        .QN(n15502) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n1540), .CK(CK), .RN(n14605), .Q(n3685), 
        .QN(n15503) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n1249), .CK(CK), .RN(n14607), .Q(n9335), 
        .QN(n15817) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n1248), .CK(CK), .RN(n14606), .Q(n9334), 
        .QN(n15818) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n3394), .CK(CK), .RN(n14605), .Q(n3127), 
        .QN(n16132) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n3398), .CK(CK), .RN(n14607), .Q(n3116), 
        .QN(n16133) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n3399), .CK(CK), .RN(n14606), .Q(n3113), 
        .QN(n16134) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n3402), .CK(CK), .RN(n14605), .Q(n3112), 
        .QN(n16135) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n3403), .CK(CK), .RN(n14607), .Q(n3140), 
        .QN(n16136) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n3405), .CK(CK), .RN(n14606), .Q(n9627), 
        .QN(n16027) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n1775), .CK(CK), .RN(n14605), .Q(n3279), 
        .QN(n15932) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n3409), .CK(CK), .RN(n14607), .Q(n3868), 
        .QN(n16028) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n3412), .CK(CK), .RN(n14606), .Q(n9630), 
        .QN(n16029) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n3413), .CK(CK), .RN(n14605), .Q(n3111), 
        .QN(n16137) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n3414), .CK(CK), .RN(n14607), .Q(n9629), 
        .QN(n16030) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n3418), .CK(CK), .RN(n14606), .Q(n3098), 
        .QN(n16138) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n1917), .CK(CK), .RN(n14605), .Q(n3884), 
        .QN(n16016) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n1916), .CK(CK), .RN(n14607), .Q(n3881), 
        .QN(n16017) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n1900), .CK(CK), .RN(n14606), .Q(n3820), 
        .QN(n16021) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n1898), .CK(CK), .RN(n14605), .Q(n3946), 
        .QN(n15925) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n1897), .CK(CK), .RN(n14607), .Q(n3941), 
        .QN(n15926) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n1892), .CK(CK), .RN(n14606), .Q(n3856), 
        .QN(n16023) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n3566), .CK(CK), .RN(n14605), .Q(n3801), 
        .QN(n16076) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n3567), .CK(CK), .RN(n14607), .Q(n3799), 
        .QN(n16077) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n3571), .CK(CK), .RN(n14606), .Q(n3664), 
        .QN(n16081) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n3572), .CK(CK), .RN(n14605), .Q(n3947), 
        .QN(n15935) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n3573), .CK(CK), .RN(n14607), .Q(n3943), 
        .QN(n15936) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n3574), .CK(CK), .RN(n14606), .Q(n3380), 
        .QN(n16083) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3435), .CK(CK), .RN(n14605), .Q(n3851), 
        .QN(n15976) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3436), .CK(CK), .RN(n14607), .Q(n3638), 
        .QN(n15978) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3438), .CK(CK), .RN(n14606), .Q(n3634), 
        .QN(n15979) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n1419), .CK(CK), .RN(n14605), .Q(n3260), 
        .QN(n16257) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3589), .CK(CK), .RN(n14607), .Q(n9754), 
        .QN(n15854) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n1155), .CK(CK), .RN(n14606), .Q(n9803), 
        .QN(n15714) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n1911), .CK(CK), .RN(n14605), .Q(n3062), 
        .QN(n16062) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n1910), .CK(CK), .RN(n14607), .Q(n9466), 
        .QN(n16063) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n1904), .CK(CK), .RN(n14606), .Q(n3957), 
        .QN(n15943) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n1902), .CK(CK), .RN(n14605), .Q(n3061), 
        .QN(n16065) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n1901), .CK(CK), .RN(n14607), .Q(n3060), 
        .QN(n16066) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n1899), .CK(CK), .RN(n14606), .Q(n3948), 
        .QN(n15944) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n1896), .CK(CK), .RN(n14605), .Q(n3231), 
        .QN(n15945) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n1894), .CK(CK), .RN(n14607), .Q(n3212), 
        .QN(n15947) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n1680), .CK(CK), .RN(n14606), .Q(n3955), 
        .QN(n15931) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n1558), .CK(CK), .RN(n14605), .Q(n9546), 
        .QN(n15585) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n1456), .CK(CK), .RN(n14607), .Q(n3828), 
        .QN(n15798) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n1451), .CK(CK), .RN(n14606), .Q(n3827), 
        .QN(n15806) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n1747), .CK(CK), .RN(n14605), .Q(n9759), 
        .QN(n15842) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n1743), .CK(CK), .RN(n14607), .Q(n9336), 
        .QN(n15865) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n1593), .CK(CK), .RN(n14606), .Q(n3635), 
        .QN(n15748) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n1586), .CK(CK), .RN(n14605), .Q(n3650), 
        .QN(n15749) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3584), .CK(CK), .RN(n14607), .Q(n9646), 
        .QN(n16266) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3585), .CK(CK), .RN(n14606), .Q(n9645), 
        .QN(n16267) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n1887), .CK(CK), .RN(n14605), .Q(n3305), 
        .QN(n16039) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n1625), .CK(CK), .RN(n14607), .Q(n3313), 
        .QN(n15539) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n1619), .CK(CK), .RN(n14606), .Q(n3083), 
        .QN(n15628) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n1618), .CK(CK), .RN(n14605), .Q(n3287), 
        .QN(n15540) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n1514), .CK(CK), .RN(n14607), .Q(n9766), 
        .QN(n15765) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n1513), .CK(CK), .RN(n14606), .Q(n9767), 
        .QN(n15766) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n1577), .CK(CK), .RN(n14605), .Q(n3131), 
        .QN(n15731) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3444), .CK(CK), .RN(n14607), .Q(n3652), 
        .QN(n16255) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3448), .CK(CK), .RN(n14606), .Q(n3665), 
        .QN(n16256) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n1950), .CK(CK), .RN(n14605), .Q(n3924), 
        .QN(n15550) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n1946), .CK(CK), .RN(n14607), .Q(n3918), 
        .QN(n15551) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n1944), .CK(CK), .RN(n14606), .Q(n3894), 
        .QN(n15553) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n1940), .CK(CK), .RN(n14605), .Q(n3888), 
        .QN(n15554) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n1927), .CK(CK), .RN(n14607), .Q(n3790), 
        .QN(n15556) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n1922), .CK(CK), .RN(n14606), .Q(n3663), 
        .QN(n15557) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3514), .CK(CK), .RN(n14605), .Q(n3639), 
        .QN(n16106) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3515), .CK(CK), .RN(n14607), .Q(n3292), 
        .QN(n16107) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3516), .CK(CK), .RN(n14606), .Q(n3291), 
        .QN(n16108) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3518), .CK(CK), .RN(n14605), .Q(n3290), 
        .QN(n16111) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3519), .CK(CK), .RN(n14607), .Q(n9664), 
        .QN(n16113) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3521), .CK(CK), .RN(n14606), .Q(n3289), 
        .QN(n16114) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3524), .CK(CK), .RN(n14605), .Q(n3637), 
        .QN(n16115) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3525), .CK(CK), .RN(n14607), .Q(n3296), 
        .QN(n16042) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3530), .CK(CK), .RN(n14606), .Q(n3689), 
        .QN(n16117) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3531), .CK(CK), .RN(n14605), .Q(n3808), 
        .QN(n16118) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n1859), .CK(CK), .RN(n14607), .Q(n3688), 
        .QN(n16045) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n1823), .CK(CK), .RN(n14606), .Q(n3865), 
        .QN(n15564) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n1537), .CK(CK), .RN(n14605), .Q(n3815), 
        .QN(n15754) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n1536), .CK(CK), .RN(n14607), .Q(n3837), 
        .QN(n15755) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n1943), .CK(CK), .RN(n14606), .Q(n3875), 
        .QN(n15743) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n1934), .CK(CK), .RN(n14605), .Q(n3298), 
        .QN(n15744) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n1933), .CK(CK), .RN(n14607), .Q(n3286), 
        .QN(n15745) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n1409), .CK(CK), .RN(n14606), .Q(n3974), 
        .QN(n15439) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n1408), .CK(CK), .RN(n14605), .Q(n3973), 
        .QN(n15440) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3420), .CK(CK), .RN(n14607), .Q(n9788), 
        .QN(n16200) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3421), .CK(CK), .RN(n14606), .Q(n9787), 
        .QN(n16201) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3422), .CK(CK), .RN(n14605), .Q(n9786), 
        .QN(n16202) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3423), .CK(CK), .RN(n14607), .Q(n9785), 
        .QN(n16203) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3427), .CK(CK), .RN(n14606), .Q(n9784), 
        .QN(n16204) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3430), .CK(CK), .RN(n14605), .Q(n9783), 
        .QN(n16205) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n1552), .CK(CK), .RN(n14607), .Q(n9563), 
        .QN(n15582) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n1951), .CK(CK), .RN(n14606), .Q(n9473), 
        .QN(n15742) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n1825), .CK(CK), .RN(n14605), .Q(n3645), 
        .QN(n15533) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n1824), .CK(CK), .RN(n14607), .Q(n3869), 
        .QN(n15534) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n1814), .CK(CK), .RN(n14606), .Q(n3789), 
        .QN(n15638) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n3392), .CK(CK), .RN(n14605), .Q(n3144), 
        .QN(n16033) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n3393), .CK(CK), .RN(n14607), .Q(n3143), 
        .QN(n16034) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n1630), .CK(CK), .RN(n14606), .Q(n3706), 
        .QN(n15624) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n1626), .CK(CK), .RN(n14605), .Q(n3707), 
        .QN(n15625) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n1624), .CK(CK), .RN(n14607), .Q(n3085), 
        .QN(n15626) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n1620), .CK(CK), .RN(n14606), .Q(n3084), 
        .QN(n15627) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n1607), .CK(CK), .RN(n14605), .Q(n3079), 
        .QN(n15629) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n1602), .CK(CK), .RN(n14607), .Q(n3708), 
        .QN(n15630) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n2047), .CK(CK), .RN(n14606), .Q(n3641), 
        .QN(n15892) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n2039), .CK(CK), .RN(n14605), .Q(n3182), 
        .QN(n15913) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n2038), .CK(CK), .RN(n14607), .Q(n3160), 
        .QN(n15914) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n2030), .CK(CK), .RN(n14606), .Q(n3181), 
        .QN(n15915) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n2029), .CK(CK), .RN(n14605), .Q(n3180), 
        .QN(n15916) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n2031), .CK(CK), .RN(n14607), .Q(n3700), 
        .QN(n15899) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3614), .CK(CK), .RN(n14606), .Q(n3282), 
        .QN(n16303) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n1719), .CK(CK), .RN(n14605), .Q(n9525), 
        .QN(n16191) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3606), .CK(CK), .RN(n14607), .Q(n9523), 
        .QN(n16192) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n1710), .CK(CK), .RN(n14606), .Q(n9527), 
        .QN(n16193) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n1709), .CK(CK), .RN(n14605), .Q(n9526), 
        .QN(n16194) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n3417), .CK(CK), .RN(n14607), .Q(n3202), 
        .QN(n15955) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n1206), .CK(CK), .RN(n14606), .Q(n9874), 
        .QN(n15816) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3616), .CK(CK), .RN(n14605), .Q(n3675), 
        .QN(n16188) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3617), .CK(CK), .RN(n14607), .Q(n3261), 
        .QN(n16189) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3618), .CK(CK), .RN(n14606), .Q(n3677), 
        .QN(n16190) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n1174), .CK(CK), .RN(n14605), .Q(n9765), 
        .QN(n15853) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n1791), .CK(CK), .RN(n14607), .Q(n3178), 
        .QN(n16072) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n3400), .CK(CK), .RN(n14606), .Q(n3135), 
        .QN(n16073) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n3401), .CK(CK), .RN(n14605), .Q(n9632), 
        .QN(n16025) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n3406), .CK(CK), .RN(n14607), .Q(n3824), 
        .QN(n16074) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n3407), .CK(CK), .RN(n14606), .Q(n3822), 
        .QN(n16075) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n1519), .CK(CK), .RN(n14605), .Q(n9349), 
        .QN(n15774) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n1273), .CK(CK), .RN(n14607), .Q(n9641), 
        .QN(n16031) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n1266), .CK(CK), .RN(n14606), .Q(n9640), 
        .QN(n16032) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n1215), .CK(CK), .RN(n14605), .Q(n9858), 
        .QN(n15864) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n1529), .CK(CK), .RN(n14607), .Q(n9348), 
        .QN(n15919) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n1526), .CK(CK), .RN(n14606), .Q(n9790), 
        .QN(n15833) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n1522), .CK(CK), .RN(n14605), .Q(n9350), 
        .QN(n15920) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n1520), .CK(CK), .RN(n14607), .Q(n9495), 
        .QN(n15708) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n1515), .CK(CK), .RN(n14606), .Q(n9492), 
        .QN(n15709) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n1512), .CK(CK), .RN(n14605), .Q(n9494), 
        .QN(n15710) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n1510), .CK(CK), .RN(n14607), .Q(n9493), 
        .QN(n15712) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n1399), .CK(CK), .RN(n14606), .Q(n9835), 
        .QN(n15732) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n1390), .CK(CK), .RN(n14605), .Q(n9837), 
        .QN(n15733) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n1389), .CK(CK), .RN(n14607), .Q(n9836), 
        .QN(n15734) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n1583), .CK(CK), .RN(n14606), .Q(n3101), 
        .QN(n15645) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n2053), .CK(CK), .RN(n14605), .Q(n9851), 
        .QN(n16228) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n1481), .CK(CK), .RN(n14607), .Q(n3055), 
        .QN(n15580) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n1337), .CK(CK), .RN(n14606), .Q(n3679), 
        .QN(n16175) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n1330), .CK(CK), .RN(n14605), .Q(n3262), 
        .QN(n16176) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n1327), .CK(CK), .RN(n14607), .Q(n3265), 
        .QN(n16177) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n3595), .CK(CK), .RN(n14606), .Q(n3716), 
        .QN(n16151) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n2013), .CK(CK), .RN(n14605), .Q(n9367), 
        .QN(n15873) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n2012), .CK(CK), .RN(n14607), .Q(n9372), 
        .QN(n15874) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n2011), .CK(CK), .RN(n14606), .Q(n9369), 
        .QN(n15875) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n2005), .CK(CK), .RN(n14605), .Q(n9368), 
        .QN(n15877) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n2001), .CK(CK), .RN(n14607), .Q(n9370), 
        .QN(n15880) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n1996), .CK(CK), .RN(n14606), .Q(n9371), 
        .QN(n15881) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n1995), .CK(CK), .RN(n14605), .Q(n9397), 
        .QN(n15847) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n1994), .CK(CK), .RN(n14607), .Q(n9497), 
        .QN(n15882) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n1989), .CK(CK), .RN(n14606), .Q(n9496), 
        .QN(n15884) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n1988), .CK(CK), .RN(n14605), .Q(n9366), 
        .QN(n15885) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3546), .CK(CK), .RN(n14607), .Q(n9815), 
        .QN(n15795) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n1829), .CK(CK), .RN(n14606), .Q(n9818), 
        .QN(n15840) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n1827), .CK(CK), .RN(n14605), .Q(n9817), 
        .QN(n15841) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n1736), .CK(CK), .RN(n14607), .Q(n9777), 
        .QN(n15722) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n1734), .CK(CK), .RN(n14606), .Q(n9776), 
        .QN(n15723) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n1195), .CK(CK), .RN(n14605), .Q(n9864), 
        .QN(n15845) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n1187), .CK(CK), .RN(n14607), .Q(n9863), 
        .QN(n15668) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n1179), .CK(CK), .RN(n14606), .Q(n9743), 
        .QN(n15819) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n1173), .CK(CK), .RN(n14605), .Q(n9742), 
        .QN(n15820) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n1169), .CK(CK), .RN(n14607), .Q(n9741), 
        .QN(n15821) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3419), .CK(CK), .RN(n14606), .Q(n9381), 
        .QN(n16293) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n1725), .CK(CK), .RN(n14605), .Q(n3836), 
        .QN(n16179) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n1724), .CK(CK), .RN(n14607), .Q(n3835), 
        .QN(n16180) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n1723), .CK(CK), .RN(n14606), .Q(n3834), 
        .QN(n16181) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n1717), .CK(CK), .RN(n14605), .Q(n3830), 
        .QN(n16182) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3424), .CK(CK), .RN(n14607), .Q(n9528), 
        .QN(n16172) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n1713), .CK(CK), .RN(n14606), .Q(n3829), 
        .QN(n16183) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n1708), .CK(CK), .RN(n14605), .Q(n3207), 
        .QN(n16185) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n1707), .CK(CK), .RN(n14607), .Q(n9811), 
        .QN(n16186) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n1706), .CK(CK), .RN(n14606), .Q(n3201), 
        .QN(n16294) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3426), .CK(CK), .RN(n14605), .Q(n3814), 
        .QN(n16253) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3428), .CK(CK), .RN(n14607), .Q(n3812), 
        .QN(n16254) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n1701), .CK(CK), .RN(n14606), .Q(n3810), 
        .QN(n16304) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n1700), .CK(CK), .RN(n14605), .Q(n3809), 
        .QN(n16187) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3429), .CK(CK), .RN(n14607), .Q(n3807), 
        .QN(n16305) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3611), .CK(CK), .RN(n14606), .Q(n3644), 
        .QN(n15949) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3612), .CK(CK), .RN(n14605), .Q(n3867), 
        .QN(n15950) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n1691), .CK(CK), .RN(n14607), .Q(n3796), 
        .QN(n16046) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n1685), .CK(CK), .RN(n14606), .Q(n3726), 
        .QN(n16047) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n1681), .CK(CK), .RN(n14605), .Q(n3672), 
        .QN(n16048) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n1667), .CK(CK), .RN(n14607), .Q(n3345), 
        .QN(n15960) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n1561), .CK(CK), .RN(n14606), .Q(n9861), 
        .QN(n15584) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n1554), .CK(CK), .RN(n14605), .Q(n9860), 
        .QN(n15586) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n1547), .CK(CK), .RN(n14607), .Q(n9872), 
        .QN(n15651) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n1541), .CK(CK), .RN(n14606), .Q(n9828), 
        .QN(n15583) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n1225), .CK(CK), .RN(n14605), .Q(n9781), 
        .QN(n15830) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n1879), .CK(CK), .RN(n14607), .Q(n3115), 
        .QN(n15956) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n1878), .CK(CK), .RN(n14606), .Q(n3123), 
        .QN(n15957) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n1870), .CK(CK), .RN(n14605), .Q(n3110), 
        .QN(n15958) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n1869), .CK(CK), .RN(n14607), .Q(n3114), 
        .QN(n15959) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n1623), .CK(CK), .RN(n14606), .Q(n3960), 
        .QN(n15435) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n1622), .CK(CK), .RN(n14605), .Q(n3089), 
        .QN(n15780) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n1614), .CK(CK), .RN(n14607), .Q(n3959), 
        .QN(n15436) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n1613), .CK(CK), .RN(n14606), .Q(n3958), 
        .QN(n15437) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n1559), .CK(CK), .RN(n14605), .Q(n3892), 
        .QN(n15511) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n1550), .CK(CK), .RN(n14607), .Q(n3953), 
        .QN(n15512) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n1549), .CK(CK), .RN(n14606), .Q(n3952), 
        .QN(n15513) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n1729), .CK(CK), .RN(n14605), .Q(n9357), 
        .QN(n16291) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n1728), .CK(CK), .RN(n14607), .Q(n9356), 
        .QN(n16292) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n1459), .CK(CK), .RN(n14606), .Q(n9417), 
        .QN(n15700) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n1247), .CK(CK), .RN(n14605), .Q(n3805), 
        .QN(n15850) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3741), .CK(CK), .RN(n14607), .Q(n3909), 
        .QN(n15768) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n2051), .CK(CK), .RN(n14606), .Q(n9421), 
        .QN(n16229) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n1967), .CK(CK), .RN(n14605), .Q(n9826), 
        .QN(n15860) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n1502), .CK(CK), .RN(n14607), .Q(n9672), 
        .QN(n15678) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n1498), .CK(CK), .RN(n14606), .Q(n9673), 
        .QN(n15679) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n1496), .CK(CK), .RN(n14605), .Q(n9668), 
        .QN(n15680) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n1492), .CK(CK), .RN(n14607), .Q(n9667), 
        .QN(n15681) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n1488), .CK(CK), .RN(n14606), .Q(n3169), 
        .QN(n15504) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n1487), .CK(CK), .RN(n14605), .Q(n3975), 
        .QN(n15432) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n1479), .CK(CK), .RN(n14607), .Q(n9669), 
        .QN(n15682) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n1474), .CK(CK), .RN(n14606), .Q(n9671), 
        .QN(n15684) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3730), .CK(CK), .RN(n14605), .Q(n3903), 
        .QN(n15699) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n1343), .CK(CK), .RN(n14607), .Q(n3266), 
        .QN(n16174) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n1331), .CK(CK), .RN(n14606), .Q(n3263), 
        .QN(n16167) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n1235), .CK(CK), .RN(n14605), .Q(n9389), 
        .QN(n15909) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n3496), .CK(CK), .RN(n14607), .Q(n3331), 
        .QN(n16000) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n3497), .CK(CK), .RN(n14606), .Q(n3319), 
        .QN(n16001) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n3498), .CK(CK), .RN(n14605), .Q(n3317), 
        .QN(n16002) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n3500), .CK(CK), .RN(n14607), .Q(n3306), 
        .QN(n16003) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n3503), .CK(CK), .RN(n14606), .Q(n3281), 
        .QN(n16004) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n3505), .CK(CK), .RN(n14605), .Q(n3276), 
        .QN(n16006) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n3390), .CK(CK), .RN(n14607), .Q(n3268), 
        .QN(n16128) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n3506), .CK(CK), .RN(n14606), .Q(n3241), 
        .QN(n16052) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n3509), .CK(CK), .RN(n14605), .Q(n3238), 
        .QN(n16170) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n3510), .CK(CK), .RN(n14607), .Q(n3211), 
        .QN(n16007) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n3511), .CK(CK), .RN(n14606), .Q(n3237), 
        .QN(n16171) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n1968), .CK(CK), .RN(n14605), .Q(n9878), 
        .QN(n15715) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n1320), .CK(CK), .RN(n14607), .Q(n3217), 
        .QN(n16085) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n1318), .CK(CK), .RN(n14606), .Q(n3216), 
        .QN(n16086) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n3473), .CK(CK), .RN(n14605), .Q(n3676), 
        .QN(n16237) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n3476), .CK(CK), .RN(n14607), .Q(n3312), 
        .QN(n16238) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n3477), .CK(CK), .RN(n14606), .Q(n3678), 
        .QN(n16239) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n1919), .CK(CK), .RN(n14605), .Q(n3339), 
        .QN(n15937) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n1918), .CK(CK), .RN(n14607), .Q(n3092), 
        .QN(n15938) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n1914), .CK(CK), .RN(n14606), .Q(n3087), 
        .QN(n15939) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n1912), .CK(CK), .RN(n14605), .Q(n3086), 
        .QN(n15940) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n1908), .CK(CK), .RN(n14607), .Q(n3082), 
        .QN(n15941) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n1907), .CK(CK), .RN(n14606), .Q(n3302), 
        .QN(n15942) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n1895), .CK(CK), .RN(n14605), .Q(n3081), 
        .QN(n15946) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n1890), .CK(CK), .RN(n14607), .Q(n3080), 
        .QN(n15948) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n1903), .CK(CK), .RN(n14606), .Q(n9462), 
        .QN(n16163) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n2103), .CK(CK), .RN(n14605), .Q(n3309), 
        .QN(n15990) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n2102), .CK(CK), .RN(n14607), .Q(n3307), 
        .QN(n15991) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n2094), .CK(CK), .RN(n14606), .Q(n3278), 
        .QN(n15992) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n2093), .CK(CK), .RN(n14605), .Q(n3277), 
        .QN(n15993) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n1335), .CK(CK), .RN(n14607), .Q(n3721), 
        .QN(n16215) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3607), .CK(CK), .RN(n14606), .Q(n3723), 
        .QN(n16216) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n1326), .CK(CK), .RN(n14605), .Q(n3259), 
        .QN(n16217) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n1325), .CK(CK), .RN(n14607), .Q(n3722), 
        .QN(n16218) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n2081), .CK(CK), .RN(n14606), .Q(n9556), 
        .QN(n16234) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n2080), .CK(CK), .RN(n14605), .Q(n9555), 
        .QN(n16235) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n1642), .CK(CK), .RN(n14607), .Q(n3102), 
        .QN(n16008) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n1641), .CK(CK), .RN(n14606), .Q(n3100), 
        .QN(n16009) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n1503), .CK(CK), .RN(n14605), .Q(n9670), 
        .QN(n15677) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n1497), .CK(CK), .RN(n14607), .Q(n3971), 
        .QN(n15433) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n1490), .CK(CK), .RN(n14606), .Q(n3972), 
        .QN(n15434) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n3599), .CK(CK), .RN(n14605), .Q(n3283), 
        .QN(n16087) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n2067), .CK(CK), .RN(n14607), .Q(n9560), 
        .QN(n16101) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n2056), .CK(CK), .RN(n14606), .Q(n9559), 
        .QN(n16102) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n2054), .CK(CK), .RN(n14605), .Q(n9558), 
        .QN(n16103) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n3501), .CK(CK), .RN(n14607), .Q(n9681), 
        .QN(n16168) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n3507), .CK(CK), .RN(n14606), .Q(n3321), 
        .QN(n16169) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n3597), .CK(CK), .RN(n14605), .Q(n3285), 
        .QN(n16152) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n3598), .CK(CK), .RN(n14607), .Q(n3284), 
        .QN(n16153) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n2058), .CK(CK), .RN(n14606), .Q(n9853), 
        .QN(n16149) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n2057), .CK(CK), .RN(n14605), .Q(n9852), 
        .QN(n16150) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n1491), .CK(CK), .RN(n14607), .Q(n3172), 
        .QN(n15509) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n2079), .CK(CK), .RN(n14606), .Q(n9873), 
        .QN(n16269) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n1985), .CK(CK), .RN(n14605), .Q(n9880), 
        .QN(n15697) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n1984), .CK(CK), .RN(n14607), .Q(n9879), 
        .QN(n15698) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n1505), .CK(CK), .RN(n14606), .Q(n3134), 
        .QN(n15497) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n1504), .CK(CK), .RN(n14605), .Q(n3196), 
        .QN(n15498) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n1501), .CK(CK), .RN(n14607), .Q(n3191), 
        .QN(n15514) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n1500), .CK(CK), .RN(n14606), .Q(n3186), 
        .QN(n15515) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n1499), .CK(CK), .RN(n14605), .Q(n3176), 
        .QN(n15516) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n1493), .CK(CK), .RN(n14607), .Q(n3173), 
        .QN(n15517) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n1489), .CK(CK), .RN(n14606), .Q(n3170), 
        .QN(n15518) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n1484), .CK(CK), .RN(n14605), .Q(n3152), 
        .QN(n15519) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n1483), .CK(CK), .RN(n14607), .Q(n3151), 
        .QN(n15505) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n1477), .CK(CK), .RN(n14606), .Q(n3970), 
        .QN(n15426) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n1476), .CK(CK), .RN(n14605), .Q(n3167), 
        .QN(n15683) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n1475), .CK(CK), .RN(n14607), .Q(n3124), 
        .QN(n15531) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3463), .CK(CK), .RN(n14606), .Q(n9683), 
        .QN(n16178) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n3596), .CK(CK), .RN(n14605), .Q(n3673), 
        .QN(n16104) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n1993), .CK(CK), .RN(n14607), .Q(n9470), 
        .QN(n15883) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n1855), .CK(CK), .RN(n14606), .Q(n9825), 
        .QN(n15837) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3539), .CK(CK), .RN(n14605), .Q(n9871), 
        .QN(n15796) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3544), .CK(CK), .RN(n14607), .Q(n9870), 
        .QN(n15797) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3547), .CK(CK), .RN(n14606), .Q(n9854), 
        .QN(n15813) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n1753), .CK(CK), .RN(n14605), .Q(n9362), 
        .QN(n15718) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n1746), .CK(CK), .RN(n14607), .Q(n9363), 
        .QN(n15719) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n1599), .CK(CK), .RN(n14606), .Q(n3967), 
        .QN(n15438) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n1597), .CK(CK), .RN(n14605), .Q(n3192), 
        .QN(n15567) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n1596), .CK(CK), .RN(n14607), .Q(n3187), 
        .QN(n15568) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n1595), .CK(CK), .RN(n14606), .Q(n3177), 
        .QN(n15569) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n1589), .CK(CK), .RN(n14605), .Q(n3174), 
        .QN(n15570) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n1587), .CK(CK), .RN(n14607), .Q(n3088), 
        .QN(n15604) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n1585), .CK(CK), .RN(n14606), .Q(n3171), 
        .QN(n15571) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n1580), .CK(CK), .RN(n14605), .Q(n3168), 
        .QN(n15572) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n1579), .CK(CK), .RN(n14607), .Q(n3094), 
        .QN(n15631) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n1578), .CK(CK), .RN(n14606), .Q(n3150), 
        .QN(n15536) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n1576), .CK(CK), .RN(n14605), .Q(n3704), 
        .QN(n15675) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n1574), .CK(CK), .RN(n14607), .Q(n3713), 
        .QN(n15676) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n1573), .CK(CK), .RN(n14606), .Q(n3126), 
        .QN(n15573) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n1572), .CK(CK), .RN(n14605), .Q(n3125), 
        .QN(n15574) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n1571), .CK(CK), .RN(n14607), .Q(n3962), 
        .QN(n15455) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n1411), .CK(CK), .RN(n14606), .Q(n9647), 
        .QN(n16295) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n1214), .CK(CK), .RN(n14605), .Q(n9846), 
        .QN(n15867) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n1210), .CK(CK), .RN(n14607), .Q(n9844), 
        .QN(n15868) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n1208), .CK(CK), .RN(n14606), .Q(n9845), 
        .QN(n15869) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n1204), .CK(CK), .RN(n14605), .Q(n9843), 
        .QN(n15870) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n1191), .CK(CK), .RN(n14607), .Q(n9842), 
        .QN(n15871) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n1186), .CK(CK), .RN(n14606), .Q(n9841), 
        .QN(n15872) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3583), .CK(CK), .RN(n14605), .Q(n9481), 
        .QN(n15786) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n1598), .CK(CK), .RN(n14607), .Q(n3122), 
        .QN(n15600) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n1594), .CK(CK), .RN(n14606), .Q(n3121), 
        .QN(n15601) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n1592), .CK(CK), .RN(n14605), .Q(n3120), 
        .QN(n15602) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n1588), .CK(CK), .RN(n14607), .Q(n3119), 
        .QN(n15603) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n1575), .CK(CK), .RN(n14606), .Q(n3118), 
        .QN(n15605) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n1570), .CK(CK), .RN(n14605), .Q(n3117), 
        .QN(n15606) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n1430), .CK(CK), .RN(n14607), .Q(n3269), 
        .QN(n16308) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3449), .CK(CK), .RN(n14606), .Q(n3256), 
        .QN(n16173) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n2017), .CK(CK), .RN(n14605), .Q(n9365), 
        .QN(n15906) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n2016), .CK(CK), .RN(n14607), .Q(n9364), 
        .QN(n15907) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n1992), .CK(CK), .RN(n14606), .Q(n9399), 
        .QN(n15848) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n1990), .CK(CK), .RN(n14605), .Q(n9396), 
        .QN(n15849) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3550), .CK(CK), .RN(n14607), .Q(n9814), 
        .QN(n15716) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3552), .CK(CK), .RN(n14606), .Q(n9813), 
        .QN(n15717) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3442), .CK(CK), .RN(n14605), .Q(n3230), 
        .QN(n16208) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3615), .CK(CK), .RN(n14607), .Q(n3215), 
        .QN(n16209) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3619), .CK(CK), .RN(n14606), .Q(n3214), 
        .QN(n16211) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3620), .CK(CK), .RN(n14605), .Q(n3213), 
        .QN(n16214) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n1759), .CK(CK), .RN(n14607), .Q(n9775), 
        .QN(n15650) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n1757), .CK(CK), .RN(n14606), .Q(n9750), 
        .QN(n15652) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n1756), .CK(CK), .RN(n14605), .Q(n9748), 
        .QN(n15653) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n1755), .CK(CK), .RN(n14607), .Q(n9749), 
        .QN(n15654) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n1749), .CK(CK), .RN(n14606), .Q(n9747), 
        .QN(n15655) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n1745), .CK(CK), .RN(n14605), .Q(n9746), 
        .QN(n15656) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n1744), .CK(CK), .RN(n14607), .Q(n9779), 
        .QN(n15720) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n1740), .CK(CK), .RN(n14606), .Q(n9751), 
        .QN(n15657) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n1739), .CK(CK), .RN(n14605), .Q(n9778), 
        .QN(n15721) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n1732), .CK(CK), .RN(n14607), .Q(n9745), 
        .QN(n15658) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n1731), .CK(CK), .RN(n14606), .Q(n9500), 
        .QN(n15866) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n1584), .CK(CK), .RN(n14605), .Q(n3714), 
        .QN(n15674) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n1750), .CK(CK), .RN(n14607), .Q(n9524), 
        .QN(n15690) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n1971), .CK(CK), .RN(n14606), .Q(n9411), 
        .QN(n15834) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3455), .CK(CK), .RN(n14605), .Q(n3649), 
        .QN(n15986) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3456), .CK(CK), .RN(n14607), .Q(n3873), 
        .QN(n15987) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3464), .CK(CK), .RN(n14606), .Q(n3944), 
        .QN(n15981) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n3391), .CK(CK), .RN(n14605), .Q(n3264), 
        .QN(n15984) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n3508), .CK(CK), .RN(n14607), .Q(n3219), 
        .QN(n15985) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n1328), .CK(CK), .RN(n14606), .Q(n3218), 
        .QN(n16084) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n1323), .CK(CK), .RN(n14605), .Q(n3220), 
        .QN(n16059) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n3627), .CK(CK), .RN(n14607), .Q(n3109), 
        .QN(n15988) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n3559), .CK(CK), .RN(n14606), .Q(n3108), 
        .QN(n15989) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n3560), .CK(CK), .RN(n14605), .Q(n3099), 
        .QN(n15994) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n2009), .CK(CK), .RN(n14607), .Q(n9398), 
        .QN(n15876) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n2002), .CK(CK), .RN(n14606), .Q(n9402), 
        .QN(n15879) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n1999), .CK(CK), .RN(n14605), .Q(n9401), 
        .QN(n15822) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3534), .CK(CK), .RN(n14607), .Q(n9824), 
        .QN(n15809) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3538), .CK(CK), .RN(n14606), .Q(n9823), 
        .QN(n15810) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3540), .CK(CK), .RN(n14605), .Q(n9822), 
        .QN(n15811) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3542), .CK(CK), .RN(n14607), .Q(n9821), 
        .QN(n15812) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3551), .CK(CK), .RN(n14606), .Q(n9819), 
        .QN(n15814) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3554), .CK(CK), .RN(n14605), .Q(n9816), 
        .QN(n15815) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n1601), .CK(CK), .RN(n14607), .Q(n3149), 
        .QN(n15598) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n1600), .CK(CK), .RN(n14606), .Q(n3148), 
        .QN(n15599) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3441), .CK(CK), .RN(n14605), .Q(n3710), 
        .QN(n16297) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3443), .CK(CK), .RN(n14607), .Q(n3235), 
        .QN(n16298) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3445), .CK(CK), .RN(n14606), .Q(n3234), 
        .QN(n16299) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3446), .CK(CK), .RN(n14605), .Q(n3233), 
        .QN(n16300) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3450), .CK(CK), .RN(n14607), .Q(n3267), 
        .QN(n16270) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3452), .CK(CK), .RN(n14606), .Q(n3232), 
        .QN(n16301) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3586), .CK(CK), .RN(n14605), .Q(n9644), 
        .QN(n16219) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3454), .CK(CK), .RN(n14607), .Q(n3712), 
        .QN(n16302) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n1199), .CK(CK), .RN(n14606), .Q(n9562), 
        .QN(n15799) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3582), .CK(CK), .RN(n14605), .Q(n9483), 
        .QN(n15772) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3487), .CK(CK), .RN(n14607), .Q(n9482), 
        .QN(n15773) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3447), .CK(CK), .RN(n14606), .Q(n3223), 
        .QN(n16210) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3451), .CK(CK), .RN(n14605), .Q(n3222), 
        .QN(n16212) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3453), .CK(CK), .RN(n14607), .Q(n3221), 
        .QN(n16213) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n3469), .CK(CK), .RN(n14606), .Q(n3293), 
        .QN(n16236) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n2075), .CK(CK), .RN(n14605), .Q(n9420), 
        .QN(n16129) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n2069), .CK(CK), .RN(n14607), .Q(n9419), 
        .QN(n16130) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n2065), .CK(CK), .RN(n14606), .Q(n9418), 
        .QN(n16131) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3575), .CK(CK), .RN(n14605), .Q(n9649), 
        .QN(n16157) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3576), .CK(CK), .RN(n14607), .Q(n9651), 
        .QN(n16158) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3577), .CK(CK), .RN(n14606), .Q(n9648), 
        .QN(n16159) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3578), .CK(CK), .RN(n14605), .Q(n9652), 
        .QN(n16160) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3579), .CK(CK), .RN(n14607), .Q(n9653), 
        .QN(n16161) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3580), .CK(CK), .RN(n14606), .Q(n9650), 
        .QN(n16162) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n3467), .CK(CK), .RN(n14605), .Q(n3325), 
        .QN(n16258) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n3468), .CK(CK), .RN(n14607), .Q(n3324), 
        .QN(n16259) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n2003), .CK(CK), .RN(n14606), .Q(n9768), 
        .QN(n15878) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n1761), .CK(CK), .RN(n14605), .Q(n9394), 
        .QN(n15691) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n1760), .CK(CK), .RN(n14607), .Q(n9393), 
        .QN(n15692) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n1758), .CK(CK), .RN(n14606), .Q(n9774), 
        .QN(n15800) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n1754), .CK(CK), .RN(n14605), .Q(n9773), 
        .QN(n15801) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n1752), .CK(CK), .RN(n14607), .Q(n9772), 
        .QN(n15802) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n1748), .CK(CK), .RN(n14606), .Q(n9771), 
        .QN(n15803) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n1735), .CK(CK), .RN(n14605), .Q(n9770), 
        .QN(n15804) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n1730), .CK(CK), .RN(n14607), .Q(n9769), 
        .QN(n15805) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3613), .CK(CK), .RN(n14606), .Q(n3322), 
        .QN(n16245) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3440), .CK(CK), .RN(n14605), .Q(n3323), 
        .QN(n16246) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n1183), .CK(CK), .RN(n14607), .Q(n9498), 
        .QN(n15911) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n2000), .CK(CK), .RN(n14606), .Q(n9400), 
        .QN(n15846) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3543), .CK(CK), .RN(n14605), .Q(n9827), 
        .QN(n15838) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n1834), .CK(CK), .RN(n14607), .Q(n9820), 
        .QN(n15839) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n1431), .CK(CK), .RN(n14606), .Q(n3257), 
        .QN(n16307) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n1422), .CK(CK), .RN(n14605), .Q(n3255), 
        .QN(n16309) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n1421), .CK(CK), .RN(n14607), .Q(n3254), 
        .QN(n16310) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n1963), .CK(CK), .RN(n14606), .Q(n9866), 
        .QN(n15693) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n1960), .CK(CK), .RN(n14605), .Q(n9877), 
        .QN(n15835) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n1958), .CK(CK), .RN(n14607), .Q(n9876), 
        .QN(n15836) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n3471), .CK(CK), .RN(n14606), .Q(n9662), 
        .QN(n16230) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n3472), .CK(CK), .RN(n14605), .Q(n9661), 
        .QN(n16231) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n3592), .CK(CK), .RN(n14607), .Q(n3718), 
        .QN(n16260) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n3475), .CK(CK), .RN(n14606), .Q(n3703), 
        .QN(n16268) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n3593), .CK(CK), .RN(n14605), .Q(n3720), 
        .QN(n16261) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n3478), .CK(CK), .RN(n14607), .Q(n9660), 
        .QN(n16232) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n3481), .CK(CK), .RN(n14606), .Q(n9659), 
        .QN(n16233) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n1655), .CK(CK), .RN(n14605), .Q(n3130), 
        .QN(n16195) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n1654), .CK(CK), .RN(n14607), .Q(n3106), 
        .QN(n16196) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n1648), .CK(CK), .RN(n14606), .Q(n3069), 
        .QN(n15968) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n1646), .CK(CK), .RN(n14605), .Q(n3129), 
        .QN(n16197) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n1645), .CK(CK), .RN(n14607), .Q(n3128), 
        .QN(n16198) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n1643), .CK(CK), .RN(n14606), .Q(n3059), 
        .QN(n15969) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n1640), .CK(CK), .RN(n14605), .Q(n3058), 
        .QN(n15970) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n1638), .CK(CK), .RN(n14607), .Q(n3057), 
        .QN(n15972) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n1495), .CK(CK), .RN(n14606), .Q(n3978), 
        .QN(n15427) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n1494), .CK(CK), .RN(n14605), .Q(n3053), 
        .QN(n15632) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n1486), .CK(CK), .RN(n14607), .Q(n3977), 
        .QN(n15428) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n1485), .CK(CK), .RN(n14606), .Q(n3976), 
        .QN(n15429) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n1847), .CK(CK), .RN(n14605), .Q(n9869), 
        .QN(n15686) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n1846), .CK(CK), .RN(n14607), .Q(n9890), 
        .QN(n15687) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n1838), .CK(CK), .RN(n14606), .Q(n9868), 
        .QN(n15688) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n1837), .CK(CK), .RN(n14605), .Q(n9867), 
        .QN(n15689) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n1590), .CK(CK), .RN(n14607), .Q(n3091), 
        .QN(n15781) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n3499), .CK(CK), .RN(n14606), .Q(n3315), 
        .QN(n15982) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n3502), .CK(CK), .RN(n14605), .Q(n3288), 
        .QN(n15983) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n3504), .CK(CK), .RN(n14607), .Q(n3275), 
        .QN(n16154) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n3389), .CK(CK), .RN(n14606), .Q(n3280), 
        .QN(n16005) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n2077), .CK(CK), .RN(n14605), .Q(n9850), 
        .QN(n16240) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n2076), .CK(CK), .RN(n14607), .Q(n9849), 
        .QN(n16241) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n2060), .CK(CK), .RN(n14606), .Q(n9848), 
        .QN(n16242) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n2052), .CK(CK), .RN(n14605), .Q(n9847), 
        .QN(n16243) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n1983), .CK(CK), .RN(n14607), .Q(n9547), 
        .QN(n15790) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n1977), .CK(CK), .RN(n14606), .Q(n9857), 
        .QN(n15807) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n1970), .CK(CK), .RN(n14605), .Q(n9856), 
        .QN(n15808) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n1961), .CK(CK), .RN(n14607), .Q(n9862), 
        .QN(n15792) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n1665), .CK(CK), .RN(n14606), .Q(n9655), 
        .QN(n16155) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n1664), .CK(CK), .RN(n14605), .Q(n9656), 
        .QN(n16156) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n1283), .CK(CK), .RN(n14607), .Q(n3320), 
        .QN(n16148) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n1659), .CK(CK), .RN(n14606), .Q(n3107), 
        .QN(n15996) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n1653), .CK(CK), .RN(n14605), .Q(n3104), 
        .QN(n15997) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n1649), .CK(CK), .RN(n14607), .Q(n3105), 
        .QN(n15998) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n1637), .CK(CK), .RN(n14606), .Q(n3103), 
        .QN(n15999) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n1480), .CK(CK), .RN(n14605), .Q(n3133), 
        .QN(n15506) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n1478), .CK(CK), .RN(n14607), .Q(n3132), 
        .QN(n15507) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n3495), .CK(CK), .RN(n14606), .Q(n3246), 
        .QN(n16051) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n1981), .CK(CK), .RN(n14605), .Q(n9554), 
        .QN(n15855) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n1980), .CK(CK), .RN(n14607), .Q(n9551), 
        .QN(n15856) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n1979), .CK(CK), .RN(n14606), .Q(n9553), 
        .QN(n15857) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n1973), .CK(CK), .RN(n14605), .Q(n9550), 
        .QN(n15858) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n1969), .CK(CK), .RN(n14607), .Q(n9549), 
        .QN(n15859) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n1964), .CK(CK), .RN(n14606), .Q(n9552), 
        .QN(n15861) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n1962), .CK(CK), .RN(n14605), .Q(n9883), 
        .QN(n15791) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n1957), .CK(CK), .RN(n14607), .Q(n9882), 
        .QN(n15793) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n1956), .CK(CK), .RN(n14606), .Q(n9548), 
        .QN(n15862) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n1955), .CK(CK), .RN(n14605), .Q(n9881), 
        .QN(n15794) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n1661), .CK(CK), .RN(n14607), .Q(n9615), 
        .QN(n16097) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n1660), .CK(CK), .RN(n14606), .Q(n9614), 
        .QN(n16098) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n1644), .CK(CK), .RN(n14605), .Q(n9613), 
        .QN(n16099) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n1636), .CK(CK), .RN(n14607), .Q(n9612), 
        .QN(n16100) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n3493), .CK(CK), .RN(n14606), .Q(n9685), 
        .QN(n16049) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n3494), .CK(CK), .RN(n14605), .Q(n9684), 
        .QN(n16050) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3457), .CK(CK), .RN(n14607), .Q(n3253), 
        .QN(n16053) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3458), .CK(CK), .RN(n14606), .Q(n3252), 
        .QN(n16054) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3459), .CK(CK), .RN(n14605), .Q(n3251), 
        .QN(n16055) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3460), .CK(CK), .RN(n14607), .Q(n3250), 
        .QN(n16056) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3461), .CK(CK), .RN(n14606), .Q(n3249), 
        .QN(n16057) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3462), .CK(CK), .RN(n14605), .Q(n3248), 
        .QN(n16058) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3465), .CK(CK), .RN(n14607), .Q(n3628), 
        .QN(n16010) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3466), .CK(CK), .RN(n14606), .Q(n3247), 
        .QN(n16060) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n1315), .CK(CK), .RN(n14605), .Q(n3349), 
        .QN(n16011) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n1635), .CK(CK), .RN(n14607), .Q(n3078), 
        .QN(n15995) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n3610), .CK(CK), .RN(n14606), .Q(n3070), 
        .QN(n15962) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n3555), .CK(CK), .RN(n14605), .Q(n3077), 
        .QN(n15963) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n3556), .CK(CK), .RN(n14607), .Q(n3076), 
        .QN(n15964) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n3557), .CK(CK), .RN(n14606), .Q(n3075), 
        .QN(n15965) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n3558), .CK(CK), .RN(n14605), .Q(n3074), 
        .QN(n15966) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n1651), .CK(CK), .RN(n14607), .Q(n3073), 
        .QN(n15967) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n3561), .CK(CK), .RN(n14606), .Q(n3072), 
        .QN(n15971) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n3562), .CK(CK), .RN(n14605), .Q(n3071), 
        .QN(n15973) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n3470), .CK(CK), .RN(n14607), .Q(n9603), 
        .QN(n16271) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n3474), .CK(CK), .RN(n14606), .Q(n9599), 
        .QN(n16272) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n3621), .CK(CK), .RN(n14605), .Q(n9600), 
        .QN(n16273) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n1303), .CK(CK), .RN(n14607), .Q(n9606), 
        .QN(n16274) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n3622), .CK(CK), .RN(n14606), .Q(n9598), 
        .QN(n16275) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n3623), .CK(CK), .RN(n14605), .Q(n9608), 
        .QN(n16276) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n1294), .CK(CK), .RN(n14607), .Q(n9604), 
        .QN(n16277) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n1293), .CK(CK), .RN(n14606), .Q(n9605), 
        .QN(n16278) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n3624), .CK(CK), .RN(n14605), .Q(n9609), 
        .QN(n16279) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n3479), .CK(CK), .RN(n14607), .Q(n9601), 
        .QN(n16280) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n3480), .CK(CK), .RN(n14606), .Q(n9607), 
        .QN(n16281) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n3482), .CK(CK), .RN(n14605), .Q(n9602), 
        .QN(n16282) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n2135), .CK(CK), .RN(n14607), .QN(
        n16311) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n2134), .CK(CK), .RN(n14606), .QN(
        n16199) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n2126), .CK(CK), .RN(n14605), .QN(
        n16312) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n2125), .CK(CK), .RN(n14607), .QN(
        n16313) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n3385), .CK(CK), .RN(n14606), .QN(
        n16247) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n3386), .CK(CK), .RN(n14605), .QN(
        n16248) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n3625), .CK(CK), .RN(n14607), .Q(n9395), 
        .QN(n16263) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n3388), .CK(CK), .RN(n14606), .Q(n9479), 
        .QN(n16251) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n3609), .CK(CK), .RN(n14605), .Q(n9478), 
        .QN(n16252) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n3626), .CK(CK), .RN(n14607), .Q(n9378), 
        .QN(n16206) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n2121), .CK(CK), .RN(n14606), .Q(n3817), 
        .QN(n16306) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n2143), .CK(CK), .RN(n14605), .Q(n9388), 
        .QN(n16262) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n2141), .CK(CK), .RN(n14607), .Q(n3189), 
        .QN(n16220) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n2140), .CK(CK), .RN(n14606), .Q(n3188), 
        .QN(n16221) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n2139), .CK(CK), .RN(n14605), .Q(n3185), 
        .QN(n16222) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n2133), .CK(CK), .RN(n14607), .Q(n3184), 
        .QN(n16223) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n2129), .CK(CK), .RN(n14606), .Q(n3142), 
        .QN(n16224) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n3387), .CK(CK), .RN(n14605), .Q(n9480), 
        .QN(n16249) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n2124), .CK(CK), .RN(n14607), .Q(n3821), 
        .QN(n16225) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n3608), .CK(CK), .RN(n14606), .Q(n9760), 
        .QN(n16250) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n2117), .CK(CK), .RN(n14605), .Q(n3139), 
        .QN(n16226) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n2116), .CK(CK), .RN(n14607), .Q(n3141), 
        .QN(n16227) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n2115), .CK(CK), .RN(n14606), .Q(n9472), 
        .QN(n16207) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n2142), .CK(CK), .RN(n14605), .Q(n9387), 
        .QN(n16285) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n2138), .CK(CK), .RN(n14607), .Q(n9386), 
        .QN(n16286) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n2136), .CK(CK), .RN(n14606), .Q(n9385), 
        .QN(n16287) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n2132), .CK(CK), .RN(n14605), .Q(n9384), 
        .QN(n16288) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n2119), .CK(CK), .RN(n14607), .Q(n9383), 
        .QN(n16289) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n2114), .CK(CK), .RN(n14606), .Q(n9382), 
        .QN(n16290) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n1369), .CK(CK), .RN(n14605), .Q(n3898), 
        .QN(n15751) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n1363), .CK(CK), .RN(n14607), .Q(n3146), 
        .QN(n15607) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n1362), .CK(CK), .RN(n14606), .Q(n3900), 
        .QN(n15752) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n2145), .CK(CK), .RN(n14605), .Q(n9538), 
        .QN(n16283) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n2144), .CK(CK), .RN(n14607), .Q(n9537), 
        .QN(n16284) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n1377), .CK(CK), .RN(n14606), .Q(n3832), 
        .QN(n15537) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n1376), .CK(CK), .RN(n14605), .Q(n3939), 
        .QN(n15538) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n1373), .CK(CK), .RN(n14607), .Q(n3849), 
        .QN(n15756) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n1372), .CK(CK), .RN(n14606), .Q(n3848), 
        .QN(n15757) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n1371), .CK(CK), .RN(n14605), .Q(n3847), 
        .QN(n15758) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n1365), .CK(CK), .RN(n14607), .Q(n3845), 
        .QN(n15759) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n1361), .CK(CK), .RN(n14606), .Q(n3844), 
        .QN(n15760) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n1356), .CK(CK), .RN(n14605), .Q(n3843), 
        .QN(n15761) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n1355), .CK(CK), .RN(n14607), .Q(n3876), 
        .QN(n15576) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n1349), .CK(CK), .RN(n14606), .Q(n3840), 
        .QN(n15648) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n1348), .CK(CK), .RN(n14605), .Q(n3095), 
        .QN(n15649) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n1347), .CK(CK), .RN(n14607), .Q(n3684), 
        .QN(n15542) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n1367), .CK(CK), .RN(n14606), .Q(n3897), 
        .QN(n15782) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n1366), .CK(CK), .RN(n14605), .Q(n3846), 
        .QN(n15783) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n1358), .CK(CK), .RN(n14607), .Q(n3896), 
        .QN(n15784) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n1357), .CK(CK), .RN(n14606), .Q(n3895), 
        .QN(n15785) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n1360), .CK(CK), .RN(n14605), .Q(n3880), 
        .QN(n15575) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n1359), .CK(CK), .RN(n14607), .Q(n3877), 
        .QN(n15541) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n1353), .CK(CK), .RN(n14606), .Q(n3841), 
        .QN(n15647) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n1352), .CK(CK), .RN(n14605), .Q(n3831), 
        .QN(n15577) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n1350), .CK(CK), .RN(n14607), .Q(n3696), 
        .QN(n15578) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n1375), .CK(CK), .RN(n14606), .Q(n3850), 
        .QN(n15750) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n1374), .CK(CK), .RN(n14605), .Q(n3925), 
        .QN(n15544) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n1370), .CK(CK), .RN(n14607), .Q(n3919), 
        .QN(n15545) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n1368), .CK(CK), .RN(n14606), .Q(n3899), 
        .QN(n15546) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n1364), .CK(CK), .RN(n14605), .Q(n3889), 
        .QN(n15547) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n1351), .CK(CK), .RN(n14607), .Q(n3818), 
        .QN(n15548) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n1346), .CK(CK), .RN(n14606), .Q(n3666), 
        .QN(n15549) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n1354), .CK(CK), .RN(n14605), .Q(n3842), 
        .QN(n15646) );
  NOR3_X1 U3 ( .A1(n14887), .A2(Read_two_address[1]), .A3(n15280), .ZN(n3025)
         );
  NOR3_X1 U4 ( .A1(n14887), .A2(Read_two_address[0]), .A3(n15281), .ZN(n3037)
         );
  NOR3_X1 U5 ( .A1(n15281), .A2(n14887), .A3(n15280), .ZN(n3036) );
  NOR3_X1 U6 ( .A1(Read_two_address[0]), .A2(Read_two_address[1]), .A3(n14887), 
        .ZN(n3038) );
  NOR3_X1 U7 ( .A1(Write_address[3]), .A2(Write_address[4]), .A3(n16314), .ZN(
        n1127) );
  NOR3_X1 U8 ( .A1(n15313), .A2(Write_address[4]), .A3(n16314), .ZN(n1121) );
  NOR3_X1 U9 ( .A1(n15314), .A2(Write_address[3]), .A3(n16314), .ZN(n1118) );
  NOR3_X1 U10 ( .A1(n15314), .A2(n15313), .A3(n16314), .ZN(n1101) );
  AND2_X1 U11 ( .A1(n15302), .A2(Read_one_address[2]), .ZN(n14601) );
  AND2_X1 U12 ( .A1(n1108), .A2(n1101), .ZN(n14602) );
  AND4_X1 U13 ( .A1(n2579), .A2(n2580), .A3(n2581), .A4(n2582), .ZN(n14603) );
  INV_X2 U14 ( .A(n15279), .ZN(n14604) );
  INV_X16 U15 ( .A(n14604), .ZN(n14605) );
  INV_X16 U16 ( .A(n14604), .ZN(n14606) );
  INV_X16 U17 ( .A(n14604), .ZN(n14607) );
  INV_X1 U18 ( .A(n2405), .ZN(n15292) );
  INV_X1 U19 ( .A(n1790), .ZN(n15291) );
  INV_X1 U20 ( .A(n15055), .ZN(n15051) );
  INV_X1 U21 ( .A(n15054), .ZN(n15050) );
  INV_X1 U22 ( .A(n15256), .ZN(n15247) );
  INV_X1 U23 ( .A(n15221), .ZN(n15212) );
  INV_X1 U24 ( .A(n15256), .ZN(n15246) );
  INV_X1 U25 ( .A(n15221), .ZN(n15211) );
  INV_X1 U26 ( .A(n15207), .ZN(n15197) );
  INV_X1 U27 ( .A(n15207), .ZN(n15198) );
  INV_X1 U28 ( .A(n14791), .ZN(n14781) );
  INV_X1 U29 ( .A(n14792), .ZN(n14782) );
  INV_X1 U30 ( .A(n14755), .ZN(n14746) );
  INV_X1 U31 ( .A(n14793), .ZN(n14783) );
  INV_X1 U32 ( .A(n14757), .ZN(n14748) );
  INV_X1 U33 ( .A(n14757), .ZN(n14747) );
  NAND2_X1 U34 ( .A1(n14732), .A2(n14844), .ZN(n1790) );
  NAND2_X1 U35 ( .A1(n14755), .A2(n14844), .ZN(n2405) );
  INV_X1 U36 ( .A(n15265), .ZN(n15258) );
  INV_X1 U37 ( .A(n15143), .ZN(n15135) );
  INV_X1 U38 ( .A(n15116), .ZN(n15109) );
  INV_X1 U39 ( .A(n15143), .ZN(n15136) );
  INV_X1 U40 ( .A(n15116), .ZN(n15108) );
  INV_X1 U41 ( .A(n15068), .ZN(n15060) );
  INV_X1 U42 ( .A(n15068), .ZN(n15061) );
  INV_X1 U43 ( .A(n15125), .ZN(n15118) );
  INV_X1 U44 ( .A(n15125), .ZN(n15117) );
  INV_X1 U45 ( .A(n15152), .ZN(n15145) );
  INV_X1 U46 ( .A(n15152), .ZN(n15144) );
  INV_X1 U47 ( .A(n15134), .ZN(n15126) );
  INV_X1 U48 ( .A(n15028), .ZN(n15021) );
  INV_X1 U49 ( .A(n15107), .ZN(n15099) );
  INV_X1 U50 ( .A(n15107), .ZN(n15100) );
  INV_X1 U51 ( .A(n15134), .ZN(n15127) );
  INV_X1 U52 ( .A(n15087), .ZN(n15079) );
  INV_X1 U53 ( .A(n15087), .ZN(n15080) );
  INV_X1 U54 ( .A(n15028), .ZN(n15020) );
  INV_X1 U55 ( .A(n15008), .ZN(n15000) );
  INV_X1 U56 ( .A(n15008), .ZN(n15001) );
  INV_X1 U57 ( .A(n15265), .ZN(n15257) );
  BUF_X1 U58 ( .A(n14602), .Z(n15055) );
  BUF_X1 U59 ( .A(n14602), .Z(n15054) );
  BUF_X1 U60 ( .A(n15053), .Z(n15056) );
  BUF_X1 U61 ( .A(n14602), .Z(n15052) );
  BUF_X1 U62 ( .A(n15245), .Z(n15256) );
  BUF_X1 U63 ( .A(n15210), .Z(n15221) );
  BUF_X1 U64 ( .A(n15196), .Z(n15207) );
  BUF_X1 U65 ( .A(n14957), .Z(n14956) );
  BUF_X1 U66 ( .A(n15019), .Z(n15018) );
  BUF_X1 U67 ( .A(n14989), .Z(n14988) );
  BUF_X1 U68 ( .A(n15098), .Z(n15097) );
  BUF_X1 U69 ( .A(n15163), .Z(n15162) );
  BUF_X1 U70 ( .A(n14978), .Z(n14977) );
  BUF_X1 U71 ( .A(n15039), .Z(n15038) );
  BUF_X1 U72 ( .A(n15098), .Z(n15090) );
  BUF_X1 U73 ( .A(n15097), .Z(n15089) );
  BUF_X1 U74 ( .A(n15098), .Z(n15093) );
  BUF_X1 U75 ( .A(n15097), .Z(n15092) );
  BUF_X1 U76 ( .A(n15098), .Z(n15091) );
  BUF_X1 U77 ( .A(n15163), .Z(n15154) );
  BUF_X1 U78 ( .A(n15162), .Z(n15155) );
  BUF_X1 U79 ( .A(n15232), .Z(n15223) );
  BUF_X1 U80 ( .A(n15078), .Z(n15070) );
  BUF_X1 U81 ( .A(n15078), .Z(n15071) );
  BUF_X1 U82 ( .A(n15183), .Z(n15175) );
  BUF_X1 U83 ( .A(n15183), .Z(n15176) );
  BUF_X1 U84 ( .A(n15039), .Z(n15031) );
  BUF_X1 U85 ( .A(n15038), .Z(n15032) );
  BUF_X1 U86 ( .A(n15039), .Z(n15030) );
  BUF_X1 U87 ( .A(n15049), .Z(n15041) );
  BUF_X1 U88 ( .A(n15049), .Z(n15042) );
  BUF_X1 U89 ( .A(n15208), .Z(n15213) );
  BUF_X1 U90 ( .A(n15194), .Z(n15200) );
  BUF_X1 U91 ( .A(n15194), .Z(n15199) );
  BUF_X1 U92 ( .A(n14999), .Z(n14991) );
  BUF_X1 U93 ( .A(n15019), .Z(n15010) );
  BUF_X1 U94 ( .A(n14989), .Z(n14980) );
  BUF_X1 U95 ( .A(n15173), .Z(n15165) );
  BUF_X1 U96 ( .A(n14978), .Z(n14969) );
  BUF_X1 U97 ( .A(n15078), .Z(n15072) );
  BUF_X1 U98 ( .A(n14602), .Z(n15053) );
  BUF_X1 U99 ( .A(n15090), .Z(n15094) );
  BUF_X1 U100 ( .A(n15163), .Z(n15156) );
  BUF_X1 U101 ( .A(n15231), .Z(n15224) );
  BUF_X1 U102 ( .A(n15183), .Z(n15177) );
  BUF_X1 U103 ( .A(n15208), .Z(n15214) );
  BUF_X1 U104 ( .A(n15194), .Z(n15201) );
  BUF_X1 U105 ( .A(n15243), .Z(n15248) );
  BUF_X1 U106 ( .A(n15242), .Z(n15234) );
  BUF_X1 U107 ( .A(n15049), .Z(n15043) );
  BUF_X1 U108 ( .A(n14967), .Z(n14959) );
  BUF_X1 U109 ( .A(n15193), .Z(n15185) );
  BUF_X1 U110 ( .A(n15244), .Z(n15251) );
  BUF_X1 U111 ( .A(n15245), .Z(n15255) );
  BUF_X1 U112 ( .A(n15196), .Z(n15205) );
  BUF_X1 U113 ( .A(n15196), .Z(n15206) );
  BUF_X1 U114 ( .A(n15209), .Z(n15218) );
  BUF_X1 U115 ( .A(n15245), .Z(n15254) );
  BUF_X1 U116 ( .A(n15244), .Z(n15252) );
  BUF_X1 U117 ( .A(n15243), .Z(n15250) );
  BUF_X1 U118 ( .A(n15244), .Z(n15253) );
  BUF_X1 U119 ( .A(n15243), .Z(n15249) );
  BUF_X1 U120 ( .A(n15195), .Z(n15204) );
  BUF_X1 U121 ( .A(n15208), .Z(n15215) );
  BUF_X1 U122 ( .A(n15210), .Z(n15220) );
  BUF_X1 U123 ( .A(n15210), .Z(n15219) );
  BUF_X1 U124 ( .A(n15209), .Z(n15217) );
  BUF_X1 U125 ( .A(n15209), .Z(n15216) );
  BUF_X1 U126 ( .A(n15195), .Z(n15202) );
  BUF_X1 U127 ( .A(n15195), .Z(n15203) );
  BUF_X1 U128 ( .A(n14957), .Z(n14953) );
  BUF_X1 U129 ( .A(n14957), .Z(n14954) );
  BUF_X1 U130 ( .A(n14956), .Z(n14951) );
  BUF_X1 U131 ( .A(n14957), .Z(n14950) );
  BUF_X1 U132 ( .A(n14956), .Z(n14949) );
  BUF_X1 U133 ( .A(n14957), .Z(n14955) );
  BUF_X1 U134 ( .A(n14950), .Z(n14952) );
  BUF_X1 U135 ( .A(n14957), .Z(n14948) );
  BUF_X1 U136 ( .A(n15058), .Z(n15057) );
  BUF_X1 U137 ( .A(n14602), .Z(n15059) );
  BUF_X1 U138 ( .A(n14602), .Z(n15058) );
  BUF_X1 U139 ( .A(n15234), .Z(n15240) );
  BUF_X1 U140 ( .A(n15242), .Z(n15237) );
  BUF_X1 U141 ( .A(n15242), .Z(n15238) );
  BUF_X1 U142 ( .A(n15242), .Z(n15239) );
  BUF_X1 U143 ( .A(n15235), .Z(n15241) );
  BUF_X1 U144 ( .A(n15242), .Z(n15236) );
  BUF_X1 U145 ( .A(n15242), .Z(n15235) );
  BUF_X1 U146 ( .A(n15049), .Z(n15046) );
  BUF_X1 U147 ( .A(n15049), .Z(n15045) );
  BUF_X1 U148 ( .A(n15049), .Z(n15044) );
  BUF_X1 U149 ( .A(n15039), .Z(n15034) );
  BUF_X1 U150 ( .A(n15038), .Z(n15033) );
  BUF_X1 U151 ( .A(n15039), .Z(n15037) );
  BUF_X1 U152 ( .A(n15039), .Z(n15036) );
  BUF_X1 U153 ( .A(n15166), .Z(n15172) );
  BUF_X1 U154 ( .A(n15173), .Z(n15169) );
  BUF_X1 U155 ( .A(n15173), .Z(n15170) );
  BUF_X1 U156 ( .A(n15173), .Z(n15168) );
  BUF_X1 U157 ( .A(n15031), .Z(n15035) );
  BUF_X1 U158 ( .A(n15173), .Z(n15167) );
  BUF_X1 U159 ( .A(n15183), .Z(n15178) );
  BUF_X1 U160 ( .A(n15078), .Z(n15074) );
  BUF_X1 U161 ( .A(n15078), .Z(n15075) );
  BUF_X1 U162 ( .A(n15175), .Z(n15182) );
  BUF_X1 U163 ( .A(n15043), .Z(n15048) );
  BUF_X1 U164 ( .A(n15046), .Z(n15047) );
  BUF_X1 U165 ( .A(n15098), .Z(n15095) );
  BUF_X1 U166 ( .A(n15169), .Z(n15171) );
  BUF_X1 U167 ( .A(n15173), .Z(n15166) );
  BUF_X1 U168 ( .A(n15078), .Z(n15073) );
  BUF_X1 U169 ( .A(n15183), .Z(n15180) );
  BUF_X1 U170 ( .A(n15098), .Z(n15096) );
  BUF_X1 U171 ( .A(n14978), .Z(n14976) );
  BUF_X1 U172 ( .A(n14978), .Z(n14975) );
  BUF_X1 U173 ( .A(n14978), .Z(n14974) );
  BUF_X1 U174 ( .A(n14977), .Z(n14973) );
  BUF_X1 U175 ( .A(n14969), .Z(n14972) );
  BUF_X1 U176 ( .A(n14977), .Z(n14971) );
  BUF_X1 U177 ( .A(n14978), .Z(n14970) );
  BUF_X1 U178 ( .A(n15183), .Z(n15179) );
  BUF_X1 U179 ( .A(n15177), .Z(n15181) );
  BUF_X1 U180 ( .A(n15072), .Z(n15077) );
  BUF_X1 U181 ( .A(n15074), .Z(n15076) );
  BUF_X1 U182 ( .A(n15163), .Z(n15161) );
  BUF_X1 U183 ( .A(n15163), .Z(n15160) );
  BUF_X1 U184 ( .A(n15163), .Z(n15159) );
  BUF_X1 U185 ( .A(n15162), .Z(n15158) );
  BUF_X1 U186 ( .A(n15154), .Z(n15157) );
  BUF_X1 U187 ( .A(n15232), .Z(n15230) );
  BUF_X1 U188 ( .A(n15232), .Z(n15229) );
  BUF_X1 U189 ( .A(n15232), .Z(n15228) );
  BUF_X1 U190 ( .A(n15231), .Z(n15227) );
  BUF_X1 U191 ( .A(n15232), .Z(n15225) );
  BUF_X1 U192 ( .A(n15223), .Z(n15226) );
  BUF_X1 U193 ( .A(n15019), .Z(n15015) );
  BUF_X1 U194 ( .A(n14992), .Z(n14997) );
  BUF_X1 U195 ( .A(n15019), .Z(n15016) );
  BUF_X1 U196 ( .A(n15018), .Z(n15013) );
  BUF_X1 U197 ( .A(n15193), .Z(n15189) );
  BUF_X1 U198 ( .A(n14999), .Z(n14995) );
  BUF_X1 U199 ( .A(n14999), .Z(n14994) );
  BUF_X1 U200 ( .A(n14999), .Z(n14993) );
  BUF_X1 U201 ( .A(n15018), .Z(n15012) );
  BUF_X1 U202 ( .A(n15019), .Z(n15011) );
  BUF_X1 U203 ( .A(n15193), .Z(n15190) );
  BUF_X1 U204 ( .A(n15185), .Z(n15191) );
  BUF_X1 U205 ( .A(n15193), .Z(n15188) );
  BUF_X1 U206 ( .A(n15193), .Z(n15187) );
  BUF_X1 U207 ( .A(n14999), .Z(n14996) );
  BUF_X1 U208 ( .A(n15019), .Z(n15017) );
  BUF_X1 U209 ( .A(n15010), .Z(n15014) );
  BUF_X1 U210 ( .A(n14989), .Z(n14986) );
  BUF_X1 U211 ( .A(n14988), .Z(n14982) );
  BUF_X1 U212 ( .A(n14989), .Z(n14984) );
  BUF_X1 U213 ( .A(n14967), .Z(n14960) );
  BUF_X1 U214 ( .A(n14988), .Z(n14983) );
  BUF_X1 U215 ( .A(n15186), .Z(n15192) );
  BUF_X1 U216 ( .A(n14961), .Z(n14965) );
  BUF_X1 U217 ( .A(n14989), .Z(n14987) );
  BUF_X1 U218 ( .A(n14980), .Z(n14985) );
  BUF_X1 U219 ( .A(n14989), .Z(n14981) );
  BUF_X1 U220 ( .A(n14995), .Z(n14998) );
  BUF_X1 U221 ( .A(n14999), .Z(n14992) );
  BUF_X1 U222 ( .A(n14967), .Z(n14962) );
  BUF_X1 U223 ( .A(n14967), .Z(n14963) );
  BUF_X1 U224 ( .A(n15193), .Z(n15186) );
  BUF_X1 U225 ( .A(n14967), .Z(n14964) );
  BUF_X1 U226 ( .A(n14967), .Z(n14961) );
  BUF_X1 U227 ( .A(n14962), .Z(n14966) );
  BUF_X1 U228 ( .A(n15232), .Z(n15231) );
  NOR2_X1 U229 ( .A1(n2405), .A2(n14733), .ZN(n1860) );
  INV_X1 U230 ( .A(n14772), .ZN(n14761) );
  INV_X1 U231 ( .A(n14772), .ZN(n14762) );
  INV_X1 U232 ( .A(n14826), .ZN(n14813) );
  INV_X1 U233 ( .A(n14805), .ZN(n14797) );
  INV_X1 U234 ( .A(n14808), .ZN(n14798) );
  INV_X1 U235 ( .A(n14736), .ZN(n14731) );
  INV_X1 U236 ( .A(n14834), .ZN(n14829) );
  INV_X1 U237 ( .A(n14735), .ZN(n14729) );
  INV_X1 U238 ( .A(n14727), .ZN(n14718) );
  INV_X1 U239 ( .A(n14807), .ZN(n14799) );
  INV_X1 U240 ( .A(n14826), .ZN(n14814) );
  INV_X1 U241 ( .A(n14826), .ZN(n14811) );
  INV_X1 U242 ( .A(n14804), .ZN(n14795) );
  INV_X1 U243 ( .A(n14723), .ZN(n14717) );
  INV_X1 U244 ( .A(n14734), .ZN(n14730) );
  INV_X1 U245 ( .A(n14806), .ZN(n14796) );
  INV_X1 U246 ( .A(n14737), .ZN(n14732) );
  INV_X1 U247 ( .A(n14826), .ZN(n14816) );
  INV_X1 U248 ( .A(n2120), .ZN(n15285) );
  NAND2_X1 U249 ( .A1(n1657), .A2(n14844), .ZN(n1873) );
  INV_X1 U250 ( .A(n14769), .ZN(n14759) );
  INV_X1 U251 ( .A(n14770), .ZN(n14760) );
  INV_X1 U252 ( .A(n1650), .ZN(n15298) );
  INV_X1 U253 ( .A(n1839), .ZN(n15288) );
  INV_X1 U254 ( .A(n1835), .ZN(n15286) );
  BUF_X1 U255 ( .A(n14745), .Z(n14756) );
  BUF_X1 U256 ( .A(n14777), .Z(n14791) );
  BUF_X1 U257 ( .A(n14745), .Z(n14755) );
  BUF_X1 U258 ( .A(n14778), .Z(n14793) );
  BUF_X1 U259 ( .A(n14777), .Z(n14792) );
  BUF_X1 U260 ( .A(n14745), .Z(n14757) );
  BUF_X1 U261 ( .A(n14743), .Z(n14749) );
  BUF_X1 U262 ( .A(n14743), .Z(n14750) );
  BUF_X1 U263 ( .A(n14775), .Z(n14784) );
  BUF_X1 U264 ( .A(n14743), .Z(n14751) );
  BUF_X1 U265 ( .A(n14775), .Z(n14785) );
  BUF_X1 U266 ( .A(n14775), .Z(n14786) );
  BUF_X1 U267 ( .A(n14744), .Z(n14752) );
  BUF_X1 U268 ( .A(n14776), .Z(n14787) );
  BUF_X1 U269 ( .A(n14744), .Z(n14753) );
  BUF_X1 U270 ( .A(n14744), .Z(n14754) );
  BUF_X1 U271 ( .A(n14776), .Z(n14788) );
  BUF_X1 U272 ( .A(n14776), .Z(n14789) );
  BUF_X1 U273 ( .A(n14777), .Z(n14790) );
  INV_X1 U274 ( .A(n14826), .ZN(n14815) );
  INV_X1 U275 ( .A(n1836), .ZN(n15287) );
  INV_X1 U276 ( .A(n1788), .ZN(n15290) );
  BUF_X1 U277 ( .A(n1177), .Z(n14872) );
  BUF_X1 U278 ( .A(n1177), .Z(n14873) );
  BUF_X1 U279 ( .A(n1177), .Z(n14874) );
  INV_X1 U280 ( .A(n14849), .ZN(n14844) );
  INV_X1 U281 ( .A(n14850), .ZN(n14845) );
  BUF_X1 U282 ( .A(n1079), .Z(n15260) );
  BUF_X1 U283 ( .A(n1079), .Z(n15264) );
  BUF_X1 U284 ( .A(n1079), .Z(n15263) );
  BUF_X1 U285 ( .A(n1079), .Z(n15261) );
  BUF_X1 U286 ( .A(n1079), .Z(n15262) );
  BUF_X1 U287 ( .A(n1079), .Z(n15259) );
  BUF_X1 U288 ( .A(n14608), .Z(n15062) );
  BUF_X1 U289 ( .A(n14608), .Z(n15063) );
  BUF_X1 U290 ( .A(n14608), .Z(n15064) );
  BUF_X1 U291 ( .A(n14608), .Z(n15065) );
  BUF_X1 U292 ( .A(n14608), .Z(n15067) );
  BUF_X1 U293 ( .A(n14608), .Z(n15066) );
  BUF_X1 U294 ( .A(n14609), .Z(n15002) );
  BUF_X1 U295 ( .A(n14609), .Z(n15007) );
  BUF_X1 U296 ( .A(n14609), .Z(n15003) );
  BUF_X1 U297 ( .A(n14609), .Z(n15006) );
  BUF_X1 U298 ( .A(n14609), .Z(n15005) );
  BUF_X1 U299 ( .A(n14609), .Z(n15004) );
  BUF_X1 U300 ( .A(n14615), .Z(n15142) );
  BUF_X1 U301 ( .A(n14615), .Z(n15139) );
  BUF_X1 U302 ( .A(n14615), .Z(n15138) );
  BUF_X1 U303 ( .A(n14615), .Z(n15141) );
  BUF_X1 U304 ( .A(n14611), .Z(n15112) );
  BUF_X1 U305 ( .A(n14611), .Z(n15110) );
  BUF_X1 U306 ( .A(n14615), .Z(n15137) );
  BUF_X1 U307 ( .A(n14611), .Z(n15115) );
  BUF_X1 U308 ( .A(n14611), .Z(n15114) );
  BUF_X1 U309 ( .A(n14611), .Z(n15113) );
  BUF_X1 U310 ( .A(n14615), .Z(n15140) );
  BUF_X1 U311 ( .A(n14611), .Z(n15111) );
  BUF_X1 U312 ( .A(n14614), .Z(n15084) );
  BUF_X1 U313 ( .A(n14614), .Z(n15086) );
  BUF_X1 U314 ( .A(n14612), .Z(n15148) );
  BUF_X1 U315 ( .A(n14613), .Z(n15129) );
  BUF_X1 U316 ( .A(n14613), .Z(n15130) );
  BUF_X1 U317 ( .A(n14612), .Z(n15151) );
  BUF_X1 U318 ( .A(n14612), .Z(n15150) );
  BUF_X1 U319 ( .A(n14612), .Z(n15149) );
  BUF_X1 U320 ( .A(n14612), .Z(n15147) );
  BUF_X1 U321 ( .A(n14612), .Z(n15146) );
  BUF_X1 U322 ( .A(n14613), .Z(n15131) );
  BUF_X1 U323 ( .A(n14613), .Z(n15133) );
  BUF_X1 U324 ( .A(n14614), .Z(n15082) );
  BUF_X1 U325 ( .A(n14613), .Z(n15128) );
  BUF_X1 U326 ( .A(n14610), .Z(n15027) );
  BUF_X1 U327 ( .A(n14610), .Z(n15025) );
  BUF_X1 U328 ( .A(n14610), .Z(n15024) );
  BUF_X1 U329 ( .A(n14610), .Z(n15023) );
  BUF_X1 U330 ( .A(n14613), .Z(n15132) );
  BUF_X1 U331 ( .A(n14614), .Z(n15081) );
  BUF_X1 U332 ( .A(n14614), .Z(n15083) );
  BUF_X1 U333 ( .A(n14614), .Z(n15085) );
  BUF_X1 U334 ( .A(n14610), .Z(n15026) );
  BUF_X1 U335 ( .A(n14610), .Z(n15022) );
  BUF_X1 U336 ( .A(n14616), .Z(n15119) );
  BUF_X1 U337 ( .A(n14617), .Z(n15101) );
  BUF_X1 U338 ( .A(n14616), .Z(n15123) );
  BUF_X1 U339 ( .A(n14617), .Z(n15103) );
  BUF_X1 U340 ( .A(n14617), .Z(n15106) );
  BUF_X1 U341 ( .A(n14616), .Z(n15124) );
  BUF_X1 U342 ( .A(n14616), .Z(n15121) );
  BUF_X1 U343 ( .A(n14616), .Z(n15122) );
  BUF_X1 U344 ( .A(n14616), .Z(n15120) );
  BUF_X1 U345 ( .A(n14617), .Z(n15102) );
  BUF_X1 U346 ( .A(n14617), .Z(n15104) );
  BUF_X1 U347 ( .A(n14617), .Z(n15105) );
  BUF_X1 U348 ( .A(n1079), .Z(n15265) );
  BUF_X1 U349 ( .A(n14608), .Z(n15068) );
  BUF_X1 U350 ( .A(n14609), .Z(n15008) );
  BUF_X1 U351 ( .A(n14615), .Z(n15143) );
  BUF_X1 U352 ( .A(n14611), .Z(n15116) );
  BUF_X1 U353 ( .A(n14612), .Z(n15152) );
  BUF_X1 U354 ( .A(n14613), .Z(n15134) );
  BUF_X1 U355 ( .A(n14614), .Z(n15087) );
  BUF_X1 U356 ( .A(n14610), .Z(n15028) );
  BUF_X1 U357 ( .A(n14616), .Z(n15125) );
  BUF_X1 U358 ( .A(n14617), .Z(n15107) );
  BUF_X1 U359 ( .A(n1083), .Z(n15210) );
  BUF_X1 U360 ( .A(n1083), .Z(n15208) );
  BUF_X1 U361 ( .A(n1083), .Z(n15209) );
  BUF_X1 U362 ( .A(n1080), .Z(n15245) );
  BUF_X1 U363 ( .A(n1084), .Z(n15196) );
  BUF_X1 U364 ( .A(n1080), .Z(n15244) );
  BUF_X1 U365 ( .A(n1080), .Z(n15243) );
  BUF_X1 U366 ( .A(n1084), .Z(n15194) );
  BUF_X1 U367 ( .A(n1084), .Z(n15195) );
  INV_X1 U368 ( .A(Reset), .ZN(n15279) );
  INV_X1 U369 ( .A(n15009), .ZN(n15019) );
  INV_X1 U370 ( .A(n14979), .ZN(n14989) );
  INV_X1 U371 ( .A(n14958), .ZN(n14967) );
  INV_X1 U372 ( .A(n15233), .ZN(n15242) );
  INV_X1 U373 ( .A(n14947), .ZN(n14957) );
  INV_X1 U374 ( .A(n15040), .ZN(n15049) );
  INV_X1 U375 ( .A(n15029), .ZN(n15039) );
  INV_X1 U376 ( .A(n15174), .ZN(n15183) );
  INV_X1 U377 ( .A(n15184), .ZN(n15193) );
  INV_X1 U378 ( .A(n15069), .ZN(n15078) );
  INV_X1 U379 ( .A(n15222), .ZN(n15232) );
  INV_X1 U380 ( .A(n14968), .ZN(n14978) );
  INV_X1 U381 ( .A(n15153), .ZN(n15163) );
  INV_X1 U382 ( .A(n14990), .ZN(n14999) );
  INV_X1 U383 ( .A(n15164), .ZN(n15173) );
  INV_X1 U384 ( .A(n15088), .ZN(n15098) );
  NAND2_X1 U385 ( .A1(n2564), .A2(n14781), .ZN(n1839) );
  NAND2_X1 U386 ( .A1(n2564), .A2(n14733), .ZN(n1835) );
  NOR2_X1 U387 ( .A1(n15273), .A2(n14748), .ZN(n1657) );
  AND2_X1 U388 ( .A1(n2564), .A2(n14724), .ZN(n1771) );
  INV_X1 U389 ( .A(n1634), .ZN(n15299) );
  NAND2_X1 U390 ( .A1(n1875), .A2(n14763), .ZN(n1650) );
  INV_X1 U391 ( .A(n1875), .ZN(n15302) );
  INV_X1 U392 ( .A(n14773), .ZN(n14763) );
  BUF_X1 U393 ( .A(n14774), .Z(n14773) );
  BUF_X1 U394 ( .A(n14827), .Z(n14826) );
  NAND2_X1 U395 ( .A1(n2564), .A2(n14833), .ZN(n2120) );
  INV_X1 U396 ( .A(n1652), .ZN(n15300) );
  BUF_X1 U397 ( .A(n14773), .Z(n14769) );
  BUF_X1 U398 ( .A(n14774), .Z(n14770) );
  BUF_X1 U399 ( .A(n14601), .Z(n14735) );
  BUF_X1 U400 ( .A(n14601), .Z(n14734) );
  BUF_X1 U401 ( .A(n14601), .Z(n14736) );
  BUF_X1 U402 ( .A(n14810), .Z(n14805) );
  BUF_X1 U403 ( .A(n14810), .Z(n14804) );
  BUF_X1 U404 ( .A(n14842), .Z(n14835) );
  BUF_X1 U405 ( .A(n14841), .Z(n14834) );
  BUF_X1 U406 ( .A(n14601), .Z(n14737) );
  BUF_X1 U407 ( .A(n14721), .Z(n14724) );
  BUF_X1 U408 ( .A(n14739), .Z(n14733) );
  BUF_X1 U409 ( .A(n14843), .Z(n14836) );
  BUF_X1 U410 ( .A(n14800), .Z(n14806) );
  BUF_X1 U411 ( .A(n14728), .Z(n14723) );
  BUF_X1 U412 ( .A(n14810), .Z(n14807) );
  BUF_X1 U413 ( .A(n14843), .Z(n14837) );
  BUF_X1 U414 ( .A(n14801), .Z(n14808) );
  BUF_X1 U415 ( .A(n14728), .Z(n14725) );
  BUF_X1 U416 ( .A(n14774), .Z(n14771) );
  BUF_X1 U417 ( .A(n14773), .Z(n14772) );
  BUF_X1 U418 ( .A(n14728), .Z(n14726) );
  BUF_X1 U419 ( .A(n14601), .Z(n14742) );
  BUF_X1 U420 ( .A(n14843), .Z(n14838) );
  BUF_X1 U421 ( .A(n14840), .Z(n14833) );
  BUF_X1 U422 ( .A(n14728), .Z(n14719) );
  BUF_X1 U423 ( .A(n14728), .Z(n14720) );
  BUF_X1 U424 ( .A(n14728), .Z(n14721) );
  BUF_X1 U425 ( .A(n14720), .Z(n14722) );
  BUF_X1 U426 ( .A(n14601), .Z(n14738) );
  BUF_X1 U427 ( .A(n14601), .Z(n14739) );
  BUF_X1 U428 ( .A(n14843), .Z(n14839) );
  BUF_X1 U429 ( .A(n14843), .Z(n14840) );
  BUF_X1 U430 ( .A(n14741), .Z(n14740) );
  BUF_X1 U431 ( .A(n14728), .Z(n14727) );
  BUF_X1 U432 ( .A(n14843), .Z(n14842) );
  BUF_X1 U433 ( .A(n14601), .Z(n14741) );
  BUF_X1 U434 ( .A(n14827), .Z(n14825) );
  BUF_X1 U435 ( .A(n1663), .Z(n14743) );
  BUF_X1 U436 ( .A(n1663), .Z(n14744) );
  BUF_X1 U437 ( .A(n1663), .Z(n14745) );
  BUF_X1 U438 ( .A(n14780), .Z(n14776) );
  BUF_X1 U439 ( .A(n14779), .Z(n14777) );
  BUF_X1 U440 ( .A(n14780), .Z(n14775) );
  BUF_X1 U441 ( .A(n14779), .Z(n14778) );
  AND2_X1 U442 ( .A1(n2564), .A2(n14768), .ZN(n1793) );
  INV_X1 U443 ( .A(n15272), .ZN(n15269) );
  NAND2_X1 U444 ( .A1(n2564), .A2(n14803), .ZN(n1836) );
  AND2_X1 U445 ( .A1(n2564), .A2(n14826), .ZN(n1826) );
  INV_X1 U446 ( .A(n15274), .ZN(n15270) );
  NAND2_X1 U447 ( .A1(n15293), .A2(n15269), .ZN(n2187) );
  BUF_X1 U448 ( .A(n14810), .Z(n14809) );
  BUF_X1 U449 ( .A(n14767), .Z(n14768) );
  BUF_X1 U450 ( .A(n14839), .Z(n14832) );
  BUF_X1 U451 ( .A(n14839), .Z(n14831) );
  BUF_X1 U452 ( .A(n14839), .Z(n14830) );
  BUF_X1 U453 ( .A(n14810), .Z(n14800) );
  BUF_X1 U454 ( .A(n14774), .Z(n14764) );
  BUF_X1 U455 ( .A(n14774), .Z(n14765) );
  BUF_X1 U456 ( .A(n14774), .Z(n14766) );
  BUF_X1 U457 ( .A(n14805), .Z(n14802) );
  BUF_X1 U458 ( .A(n14810), .Z(n14801) );
  BUF_X1 U459 ( .A(n14805), .Z(n14803) );
  BUF_X1 U460 ( .A(n14774), .Z(n14767) );
  BUF_X1 U461 ( .A(n14827), .Z(n14817) );
  BUF_X1 U462 ( .A(n14827), .Z(n14818) );
  BUF_X1 U463 ( .A(n14824), .Z(n14819) );
  BUF_X1 U464 ( .A(n14827), .Z(n14822) );
  BUF_X1 U465 ( .A(n14823), .Z(n14820) );
  BUF_X1 U466 ( .A(n14818), .Z(n14823) );
  BUF_X1 U467 ( .A(n14817), .Z(n14821) );
  BUF_X1 U468 ( .A(n14843), .Z(n14841) );
  BUF_X1 U469 ( .A(n14825), .Z(n14824) );
  NAND2_X1 U470 ( .A1(n15278), .A2(n14619), .ZN(n1788) );
  BUF_X1 U471 ( .A(n1170), .Z(n14881) );
  BUF_X1 U472 ( .A(n1178), .Z(n14869) );
  BUF_X1 U473 ( .A(n1170), .Z(n14882) );
  BUF_X1 U474 ( .A(n1178), .Z(n14870) );
  BUF_X1 U475 ( .A(n1145), .Z(n14917) );
  BUF_X1 U476 ( .A(n1150), .Z(n14905) );
  BUF_X1 U477 ( .A(n1145), .Z(n14918) );
  BUF_X1 U478 ( .A(n1150), .Z(n14906) );
  BUF_X1 U479 ( .A(n1140), .Z(n14929) );
  BUF_X1 U480 ( .A(n1161), .Z(n14893) );
  BUF_X1 U481 ( .A(n1140), .Z(n14930) );
  BUF_X1 U482 ( .A(n1161), .Z(n14894) );
  BUF_X1 U483 ( .A(n1135), .Z(n14941) );
  BUF_X1 U484 ( .A(n1196), .Z(n14857) );
  BUF_X1 U485 ( .A(n1135), .Z(n14942) );
  BUF_X1 U486 ( .A(n1196), .Z(n14858) );
  BUF_X1 U487 ( .A(n1137), .Z(n14938) );
  BUF_X1 U488 ( .A(n1142), .Z(n14926) );
  BUF_X1 U489 ( .A(n1147), .Z(n14914) );
  BUF_X1 U490 ( .A(n1152), .Z(n14902) );
  BUF_X1 U491 ( .A(n1172), .Z(n14878) );
  BUF_X1 U492 ( .A(n1163), .Z(n14890) );
  BUF_X1 U493 ( .A(n1188), .Z(n14866) );
  BUF_X1 U494 ( .A(n1202), .Z(n14854) );
  BUF_X1 U495 ( .A(n1137), .Z(n14939) );
  BUF_X1 U496 ( .A(n1142), .Z(n14927) );
  BUF_X1 U497 ( .A(n1147), .Z(n14915) );
  BUF_X1 U498 ( .A(n1152), .Z(n14903) );
  BUF_X1 U499 ( .A(n1172), .Z(n14879) );
  BUF_X1 U500 ( .A(n1163), .Z(n14891) );
  BUF_X1 U501 ( .A(n1188), .Z(n14867) );
  BUF_X1 U502 ( .A(n1202), .Z(n14855) );
  BUF_X1 U503 ( .A(n1144), .Z(n14920) );
  BUF_X1 U504 ( .A(n1160), .Z(n14896) );
  BUF_X1 U505 ( .A(n1144), .Z(n14921) );
  BUF_X1 U506 ( .A(n1160), .Z(n14897) );
  BUF_X1 U507 ( .A(n1134), .Z(n14944) );
  BUF_X1 U508 ( .A(n1149), .Z(n14908) );
  BUF_X1 U509 ( .A(n1194), .Z(n14860) );
  BUF_X1 U510 ( .A(n1134), .Z(n14945) );
  BUF_X1 U511 ( .A(n1149), .Z(n14909) );
  BUF_X1 U512 ( .A(n1194), .Z(n14861) );
  BUF_X1 U513 ( .A(n1139), .Z(n14932) );
  BUF_X1 U514 ( .A(n1139), .Z(n14933) );
  BUF_X1 U515 ( .A(n1168), .Z(n14884) );
  BUF_X1 U516 ( .A(n1168), .Z(n14885) );
  BUF_X1 U517 ( .A(n1138), .Z(n14936) );
  BUF_X1 U518 ( .A(n1143), .Z(n14924) );
  BUF_X1 U519 ( .A(n1148), .Z(n14912) );
  BUF_X1 U520 ( .A(n1153), .Z(n14900) );
  BUF_X1 U521 ( .A(n1176), .Z(n14876) );
  BUF_X1 U522 ( .A(n1189), .Z(n14864) );
  BUF_X1 U523 ( .A(n1205), .Z(n14852) );
  BUF_X1 U524 ( .A(n1138), .Z(n14935) );
  BUF_X1 U525 ( .A(n1143), .Z(n14923) );
  BUF_X1 U526 ( .A(n1148), .Z(n14911) );
  BUF_X1 U527 ( .A(n1153), .Z(n14899) );
  BUF_X1 U528 ( .A(n1176), .Z(n14875) );
  BUF_X1 U529 ( .A(n1189), .Z(n14863) );
  BUF_X1 U530 ( .A(n1205), .Z(n14851) );
  BUF_X1 U531 ( .A(n1170), .Z(n14883) );
  BUF_X1 U532 ( .A(n1178), .Z(n14871) );
  BUF_X1 U533 ( .A(n1145), .Z(n14919) );
  BUF_X1 U534 ( .A(n1150), .Z(n14907) );
  BUF_X1 U535 ( .A(n1140), .Z(n14931) );
  BUF_X1 U536 ( .A(n1161), .Z(n14895) );
  BUF_X1 U537 ( .A(n1135), .Z(n14943) );
  BUF_X1 U538 ( .A(n1196), .Z(n14859) );
  BUF_X1 U539 ( .A(n1137), .Z(n14940) );
  BUF_X1 U540 ( .A(n1142), .Z(n14928) );
  BUF_X1 U541 ( .A(n1152), .Z(n14904) );
  BUF_X1 U542 ( .A(n1147), .Z(n14916) );
  BUF_X1 U543 ( .A(n1172), .Z(n14880) );
  BUF_X1 U544 ( .A(n1163), .Z(n14892) );
  BUF_X1 U545 ( .A(n1188), .Z(n14868) );
  BUF_X1 U546 ( .A(n1202), .Z(n14856) );
  BUF_X1 U547 ( .A(n1144), .Z(n14922) );
  BUF_X1 U548 ( .A(n1160), .Z(n14898) );
  BUF_X1 U549 ( .A(n1134), .Z(n14946) );
  BUF_X1 U550 ( .A(n1149), .Z(n14910) );
  BUF_X1 U551 ( .A(n1194), .Z(n14862) );
  BUF_X1 U552 ( .A(n1139), .Z(n14934) );
  BUF_X1 U553 ( .A(n1168), .Z(n14886) );
  BUF_X1 U554 ( .A(n1138), .Z(n14937) );
  BUF_X1 U555 ( .A(n1143), .Z(n14925) );
  BUF_X1 U556 ( .A(n1148), .Z(n14913) );
  BUF_X1 U557 ( .A(n1153), .Z(n14901) );
  BUF_X1 U558 ( .A(n1176), .Z(n14877) );
  BUF_X1 U559 ( .A(n1189), .Z(n14865) );
  BUF_X1 U560 ( .A(n1205), .Z(n14853) );
  NAND2_X1 U561 ( .A1(n3032), .A2(n3036), .ZN(n1177) );
  NOR3_X1 U562 ( .A1(n15311), .A2(n15304), .A3(n15312), .ZN(n1100) );
  BUF_X1 U563 ( .A(n15322), .Z(n14641) );
  BUF_X1 U564 ( .A(n15329), .Z(n14662) );
  BUF_X1 U565 ( .A(n15326), .Z(n14653) );
  BUF_X1 U566 ( .A(n15327), .Z(n14656) );
  BUF_X1 U567 ( .A(n15336), .Z(n14683) );
  BUF_X1 U568 ( .A(n15323), .Z(n14644) );
  BUF_X1 U569 ( .A(n15331), .Z(n14669) );
  BUF_X1 U570 ( .A(n15338), .Z(n14690) );
  BUF_X1 U571 ( .A(n15318), .Z(n14630) );
  BUF_X1 U572 ( .A(n15324), .Z(n14648) );
  BUF_X1 U573 ( .A(n15335), .Z(n14681) );
  BUF_X1 U574 ( .A(n15323), .Z(n14645) );
  BUF_X1 U575 ( .A(n15329), .Z(n14663) );
  BUF_X1 U576 ( .A(n15328), .Z(n14660) );
  BUF_X1 U577 ( .A(n15319), .Z(n14633) );
  BUF_X1 U578 ( .A(n15321), .Z(n14639) );
  BUF_X1 U579 ( .A(n15332), .Z(n14672) );
  BUF_X1 U580 ( .A(n15326), .Z(n14654) );
  BUF_X1 U581 ( .A(n15327), .Z(n14657) );
  BUF_X1 U582 ( .A(n15336), .Z(n14684) );
  BUF_X1 U583 ( .A(n15322), .Z(n14642) );
  BUF_X1 U584 ( .A(n15330), .Z(n14666) );
  BUF_X1 U585 ( .A(n15334), .Z(n14678) );
  BUF_X1 U586 ( .A(n15340), .Z(n14696) );
  BUF_X1 U587 ( .A(n15315), .Z(n14621) );
  BUF_X1 U588 ( .A(n15320), .Z(n14636) );
  BUF_X1 U589 ( .A(n15333), .Z(n14675) );
  BUF_X1 U590 ( .A(n15337), .Z(n14687) );
  BUF_X1 U591 ( .A(n15339), .Z(n14693) );
  BUF_X1 U592 ( .A(n15343), .Z(n14705) );
  BUF_X1 U593 ( .A(n15344), .Z(n14708) );
  BUF_X1 U594 ( .A(n15317), .Z(n14627) );
  BUF_X1 U595 ( .A(n15325), .Z(n14651) );
  BUF_X1 U596 ( .A(n15341), .Z(n14699) );
  BUF_X1 U597 ( .A(n15342), .Z(n14702) );
  BUF_X1 U598 ( .A(n15345), .Z(n14711) );
  BUF_X1 U599 ( .A(n15346), .Z(n14714) );
  BUF_X1 U600 ( .A(n1167), .Z(n14887) );
  NAND2_X1 U601 ( .A1(n1100), .A2(n1101), .ZN(n1079) );
  BUF_X1 U602 ( .A(n15316), .Z(n14623) );
  BUF_X1 U603 ( .A(n1167), .Z(n14888) );
  BUF_X1 U604 ( .A(n15344), .Z(n14707) );
  BUF_X1 U605 ( .A(n15345), .Z(n14710) );
  BUF_X1 U606 ( .A(n15346), .Z(n14713) );
  BUF_X1 U607 ( .A(n15316), .Z(n14624) );
  BUF_X1 U608 ( .A(n15318), .Z(n14629) );
  BUF_X1 U609 ( .A(n15330), .Z(n14665) );
  BUF_X1 U610 ( .A(n15334), .Z(n14677) );
  BUF_X1 U611 ( .A(n15340), .Z(n14695) );
  BUF_X1 U612 ( .A(n15317), .Z(n14626) );
  BUF_X1 U613 ( .A(n15325), .Z(n14650) );
  BUF_X1 U614 ( .A(n15341), .Z(n14698) );
  BUF_X1 U615 ( .A(n15342), .Z(n14701) );
  BUF_X1 U616 ( .A(n15315), .Z(n14620) );
  BUF_X1 U617 ( .A(n15320), .Z(n14635) );
  BUF_X1 U618 ( .A(n15333), .Z(n14674) );
  BUF_X1 U619 ( .A(n15337), .Z(n14686) );
  BUF_X1 U620 ( .A(n15339), .Z(n14692) );
  BUF_X1 U621 ( .A(n15343), .Z(n14704) );
  BUF_X1 U622 ( .A(n15328), .Z(n14659) );
  BUF_X1 U623 ( .A(n15335), .Z(n14680) );
  BUF_X1 U624 ( .A(n15331), .Z(n14668) );
  BUF_X1 U625 ( .A(n15338), .Z(n14689) );
  BUF_X1 U626 ( .A(n15324), .Z(n14647) );
  BUF_X1 U627 ( .A(n15332), .Z(n14671) );
  BUF_X1 U628 ( .A(n15319), .Z(n14632) );
  BUF_X1 U629 ( .A(n15321), .Z(n14638) );
  BUF_X1 U630 ( .A(n15316), .Z(n14625) );
  NAND2_X1 U631 ( .A1(n1109), .A2(n1101), .ZN(n1080) );
  BUF_X1 U632 ( .A(n15334), .Z(n14679) );
  BUF_X1 U633 ( .A(n15317), .Z(n14628) );
  BUF_X1 U634 ( .A(n15318), .Z(n14631) );
  BUF_X1 U635 ( .A(n15325), .Z(n14652) );
  BUF_X1 U636 ( .A(n15330), .Z(n14667) );
  BUF_X1 U637 ( .A(n15340), .Z(n14697) );
  BUF_X1 U638 ( .A(n15341), .Z(n14700) );
  BUF_X1 U639 ( .A(n15342), .Z(n14703) );
  BUF_X1 U640 ( .A(n15345), .Z(n14712) );
  BUF_X1 U641 ( .A(n15346), .Z(n14715) );
  BUF_X1 U642 ( .A(n1167), .Z(n14889) );
  BUF_X1 U643 ( .A(n15331), .Z(n14670) );
  BUF_X1 U644 ( .A(n15338), .Z(n14691) );
  NAND2_X1 U645 ( .A1(n1117), .A2(n1121), .ZN(n1083) );
  NAND2_X1 U646 ( .A1(n1114), .A2(n1127), .ZN(n1084) );
  BUF_X1 U647 ( .A(n15328), .Z(n14661) );
  BUF_X1 U648 ( .A(n15344), .Z(n14709) );
  BUF_X1 U649 ( .A(n15319), .Z(n14634) );
  BUF_X1 U650 ( .A(n15321), .Z(n14640) );
  BUF_X1 U651 ( .A(n15324), .Z(n14649) );
  BUF_X1 U652 ( .A(n15332), .Z(n14673) );
  BUF_X1 U653 ( .A(n15335), .Z(n14682) );
  BUF_X1 U654 ( .A(n15323), .Z(n14646) );
  BUF_X1 U655 ( .A(n15322), .Z(n14643) );
  BUF_X1 U656 ( .A(n14603), .Z(n14850) );
  BUF_X1 U657 ( .A(n15329), .Z(n14664) );
  BUF_X1 U658 ( .A(n15315), .Z(n14622) );
  BUF_X1 U659 ( .A(n15320), .Z(n14637) );
  BUF_X1 U660 ( .A(n15339), .Z(n14694) );
  BUF_X1 U661 ( .A(n15343), .Z(n14706) );
  BUF_X1 U662 ( .A(n15333), .Z(n14676) );
  BUF_X1 U663 ( .A(n15337), .Z(n14688) );
  BUF_X1 U664 ( .A(n15326), .Z(n14655) );
  BUF_X1 U665 ( .A(n15327), .Z(n14658) );
  BUF_X1 U666 ( .A(n15336), .Z(n14685) );
  BUF_X1 U667 ( .A(n14603), .Z(n14849) );
  BUF_X1 U668 ( .A(n14603), .Z(n14846) );
  BUF_X1 U669 ( .A(n14603), .Z(n14848) );
  BUF_X1 U670 ( .A(n14603), .Z(n14847) );
  BUF_X1 U671 ( .A(n1122), .Z(n14990) );
  NAND2_X1 U672 ( .A1(n1108), .A2(n1121), .ZN(n1122) );
  BUF_X1 U673 ( .A(n1088), .Z(n15153) );
  NAND2_X1 U674 ( .A1(n1114), .A2(n1121), .ZN(n1088) );
  BUF_X1 U675 ( .A(n1124), .Z(n14968) );
  NAND2_X1 U676 ( .A1(n1111), .A2(n1121), .ZN(n1124) );
  BUF_X1 U677 ( .A(n1082), .Z(n15222) );
  NAND2_X1 U678 ( .A1(n1113), .A2(n1118), .ZN(n1082) );
  BUF_X1 U679 ( .A(n1097), .Z(n15069) );
  NAND2_X1 U680 ( .A1(n1108), .A2(n1118), .ZN(n1097) );
  BUF_X1 U681 ( .A(n1085), .Z(n15184) );
  NAND2_X1 U682 ( .A1(n1115), .A2(n1101), .ZN(n1085) );
  BUF_X1 U683 ( .A(n1095), .Z(n15088) );
  NAND2_X1 U684 ( .A1(n1115), .A2(n1127), .ZN(n1095) );
  BUF_X1 U685 ( .A(n1087), .Z(n15164) );
  NAND2_X1 U686 ( .A1(n1113), .A2(n1127), .ZN(n1087) );
  BUF_X1 U687 ( .A(n1086), .Z(n15174) );
  NAND2_X1 U688 ( .A1(n1114), .A2(n1101), .ZN(n1086) );
  BUF_X1 U689 ( .A(n1112), .Z(n15029) );
  NAND2_X1 U690 ( .A1(n1113), .A2(n1101), .ZN(n1112) );
  BUF_X1 U691 ( .A(n1110), .Z(n15040) );
  NAND2_X1 U692 ( .A1(n1111), .A2(n1101), .ZN(n1110) );
  BUF_X1 U693 ( .A(n1119), .Z(n15009) );
  NAND2_X1 U694 ( .A1(n1118), .A2(n1109), .ZN(n1119) );
  BUF_X1 U695 ( .A(n1123), .Z(n14979) );
  NAND2_X1 U696 ( .A1(n1121), .A2(n1109), .ZN(n1123) );
  BUF_X1 U697 ( .A(n1125), .Z(n14958) );
  NAND2_X1 U698 ( .A1(n1121), .A2(n1113), .ZN(n1125) );
  BUF_X1 U699 ( .A(n1126), .Z(n14947) );
  NAND2_X1 U700 ( .A1(n1127), .A2(n1100), .ZN(n1126) );
  BUF_X1 U701 ( .A(n1081), .Z(n15233) );
  NAND2_X1 U702 ( .A1(n1127), .A2(n1109), .ZN(n1081) );
  AND2_X1 U703 ( .A1(n1118), .A2(n1100), .ZN(n14608) );
  AND2_X1 U704 ( .A1(n1121), .A2(n1100), .ZN(n14609) );
  AND2_X1 U705 ( .A1(n1117), .A2(n1101), .ZN(n14610) );
  AND2_X1 U706 ( .A1(n1114), .A2(n1118), .ZN(n14611) );
  AND2_X1 U707 ( .A1(n1117), .A2(n1118), .ZN(n14612) );
  AND2_X1 U708 ( .A1(n1115), .A2(n1118), .ZN(n14613) );
  AND2_X1 U709 ( .A1(n1111), .A2(n1118), .ZN(n14614) );
  AND2_X1 U710 ( .A1(n1115), .A2(n1121), .ZN(n14615) );
  AND2_X1 U711 ( .A1(n1108), .A2(n1127), .ZN(n14616) );
  AND2_X1 U712 ( .A1(n1111), .A2(n1127), .ZN(n14617) );
  NAND2_X1 U713 ( .A1(n15303), .A2(n15301), .ZN(n1652) );
  AOI222_X1 U714 ( .A1(n14724), .A2(n16265), .B1(n14824), .B2(n15749), .C1(
        n14742), .C2(n16176), .ZN(n2286) );
  AOI222_X1 U715 ( .A1(n14819), .A2(n15645), .B1(n14772), .B2(n15860), .C1(
        n14741), .C2(n16177), .ZN(n2339) );
  AOI222_X1 U716 ( .A1(n14768), .A2(n15508), .B1(n14727), .B2(n16095), .C1(
        n14809), .C2(n16228), .ZN(n2512) );
  AOI222_X1 U717 ( .A1(n14768), .A2(n15532), .B1(n14809), .B2(n16229), .C1(
        n14748), .C2(n15714), .ZN(n2551) );
  AOI222_X1 U718 ( .A1(n14807), .A2(n16149), .B1(n14727), .B2(n15953), .C1(
        n14825), .C2(n15669), .ZN(n2422) );
  AOI222_X1 U719 ( .A1(n14723), .A2(n16264), .B1(n14824), .B2(n15748), .C1(
        n14742), .C2(n16175), .ZN(n2157) );
  AOI222_X1 U720 ( .A1(n14837), .A2(n15671), .B1(n14726), .B2(n16038), .C1(
        n14782), .C2(n16257), .ZN(n2402) );
  OAI222_X1 U721 ( .A1(n16144), .A2(n1835), .B1(n15896), .B2(n1836), .C1(
        n15611), .C2(n1839), .ZN(n2237) );
  OAI222_X1 U722 ( .A1(n16142), .A2(n1835), .B1(n15894), .B2(n1836), .C1(
        n15609), .C2(n1839), .ZN(n2098) );
  OAI222_X1 U723 ( .A1(n16143), .A2(n1835), .B1(n15895), .B2(n1836), .C1(
        n15610), .C2(n1839), .ZN(n2161) );
  OAI222_X1 U724 ( .A1(n16146), .A2(n1835), .B1(n15902), .B2(n1836), .C1(
        n15612), .C2(n1839), .ZN(n2472) );
  OAI222_X1 U725 ( .A1(n16147), .A2(n1835), .B1(n15904), .B2(n1836), .C1(
        n15614), .C2(n1839), .ZN(n2563) );
  OAI222_X1 U726 ( .A1(n16141), .A2(n1835), .B1(n15893), .B2(n1836), .C1(
        n15608), .C2(n1839), .ZN(n1832) );
  AOI221_X1 U727 ( .B1(n2180), .B2(n2201), .C1(n2202), .C2(n2203), .A(n2204), 
        .ZN(n2200) );
  AOI211_X1 U728 ( .C1(n14747), .C2(n15853), .A(n2209), .B(n2210), .ZN(n2203)
         );
  AOI211_X1 U729 ( .C1(n14722), .C2(n15961), .A(n2211), .B(n15270), .ZN(n2202)
         );
  AOI21_X1 U730 ( .B1(n2205), .B2(n2206), .A(n2187), .ZN(n2204) );
  AOI221_X1 U731 ( .B1(n14817), .B2(n15767), .C1(n14808), .C2(n15789), .A(
        n1873), .ZN(n2506) );
  NAND2_X1 U732 ( .A1(n15347), .A2(n15303), .ZN(n1875) );
  OAI221_X1 U733 ( .B1(n14765), .B2(n15934), .C1(n15302), .C2(n15924), .A(
        n1650), .ZN(n1720) );
  OAI221_X1 U734 ( .B1(n14766), .B2(n15933), .C1(n15302), .C2(n15923), .A(
        n1650), .ZN(n1647) );
  OAI22_X1 U735 ( .A1(n15633), .A2(n1839), .B1(n15922), .B2(n1835), .ZN(n2326)
         );
  OAI22_X1 U736 ( .A1(n15613), .A2(n14784), .B1(n16140), .B2(n14730), .ZN(
        n2548) );
  OAI221_X1 U737 ( .B1(n2541), .B2(n2322), .C1(n14625), .C2(n14844), .A(n2542), 
        .ZN(N961) );
  AOI22_X1 U738 ( .A1(n2552), .A2(n2553), .B1(n2554), .B2(n2555), .ZN(n2541)
         );
  AOI221_X1 U739 ( .B1(n14737), .B2(n15542), .C1(n14781), .C2(n15531), .A(
        n2557), .ZN(n2554) );
  NAND2_X1 U740 ( .A1(n15347), .A2(n15301), .ZN(n1634) );
  AOI22_X1 U741 ( .A1(n2146), .A2(n2147), .B1(n2148), .B2(n2149), .ZN(n2137)
         );
  AOI221_X1 U742 ( .B1(n14781), .B2(n16255), .C1(n14724), .C2(n16014), .A(
        n2151), .ZN(n2147) );
  AOI211_X1 U743 ( .C1(n14767), .C2(n15552), .A(n2152), .B(n15270), .ZN(n2146)
         );
  OAI221_X1 U744 ( .B1(n15917), .B2(n14798), .C1(n16061), .C2(n14761), .A(
        n2150), .ZN(n2149) );
  AOI22_X1 U745 ( .A1(n2277), .A2(n2278), .B1(n2148), .B2(n2279), .ZN(n2276)
         );
  AOI221_X1 U746 ( .B1(n14782), .B2(n16256), .C1(n14724), .C2(n16015), .A(
        n2281), .ZN(n2278) );
  AOI211_X1 U747 ( .C1(n14768), .C2(n15555), .A(n2282), .B(n15270), .ZN(n2277)
         );
  OAI221_X1 U748 ( .B1(n15918), .B2(n14798), .C1(n16064), .C2(n14761), .A(
        n2280), .ZN(n2279) );
  AOI22_X1 U749 ( .A1(n14738), .A2(n16152), .B1(n14782), .B2(n16266), .ZN(
        n2421) );
  OAI22_X1 U750 ( .A1(n14712), .A2(n14844), .B1(n1698), .B2(n1699), .ZN(N990)
         );
  AOI221_X1 U751 ( .B1(n1726), .B2(n1727), .C1(n1737), .C2(n1762), .A(n14619), 
        .ZN(n1698) );
  AOI21_X1 U752 ( .B1(n1702), .B2(n14844), .A(n15293), .ZN(n1699) );
  AOI221_X1 U753 ( .B1(n14733), .B2(n15538), .C1(n14783), .C2(n15498), .A(
        n1763), .ZN(n1762) );
  OAI22_X1 U754 ( .A1(n14715), .A2(n14845), .B1(n1437), .B2(n1438), .ZN(N991)
         );
  AOI221_X1 U755 ( .B1(n1672), .B2(n1683), .C1(n1684), .C2(n1688), .A(n14619), 
        .ZN(n1437) );
  AOI21_X1 U756 ( .B1(n1439), .B2(n14844), .A(n15293), .ZN(n1438) );
  AOI221_X1 U757 ( .B1(n14736), .B2(n15537), .C1(n14783), .C2(n15497), .A(
        n1690), .ZN(n1688) );
  OAI22_X1 U758 ( .A1(n14679), .A2(n14845), .B1(n2216), .B2(n2217), .ZN(N979)
         );
  AOI221_X1 U759 ( .B1(n2226), .B2(n2227), .C1(n2228), .C2(n2229), .A(n14619), 
        .ZN(n2216) );
  AOI221_X1 U760 ( .B1(n2218), .B2(n2219), .C1(n2220), .C2(n2221), .A(n15293), 
        .ZN(n2217) );
  AOI221_X1 U761 ( .B1(n14735), .B2(n15759), .C1(n14783), .C2(n15517), .A(
        n2231), .ZN(n2228) );
  OAI22_X1 U762 ( .A1(n14628), .A2(n14844), .B1(n2523), .B2(n2524), .ZN(N962)
         );
  AOI221_X1 U763 ( .B1(n2533), .B2(n2534), .C1(n2535), .C2(n2536), .A(n14618), 
        .ZN(n2523) );
  AOI221_X1 U764 ( .B1(n2525), .B2(n2526), .C1(n2527), .C2(n2528), .A(n15293), 
        .ZN(n2524) );
  AOI221_X1 U765 ( .B1(n14736), .B2(n15649), .C1(n14783), .C2(n15683), .A(
        n2538), .ZN(n2535) );
  OAI22_X1 U766 ( .A1(n14631), .A2(n14845), .B1(n2504), .B2(n2505), .ZN(N963)
         );
  AOI221_X1 U767 ( .B1(n2515), .B2(n2516), .C1(n2517), .C2(n2518), .A(n14619), 
        .ZN(n2504) );
  AOI22_X1 U768 ( .A1(n2506), .A2(n2507), .B1(n2508), .B2(n14844), .ZN(n2505)
         );
  AOI221_X1 U769 ( .B1(n14737), .B2(n15648), .C1(n14783), .C2(n15426), .A(
        n2520), .ZN(n2517) );
  OAI22_X1 U770 ( .A1(n14652), .A2(n14845), .B1(n2378), .B2(n2379), .ZN(N970)
         );
  AOI221_X1 U771 ( .B1(n2388), .B2(n2389), .C1(n2390), .C2(n2391), .A(n14618), 
        .ZN(n2378) );
  AOI221_X1 U772 ( .B1(n2380), .B2(n2381), .C1(n2382), .C2(n2383), .A(n15293), 
        .ZN(n2379) );
  AOI221_X1 U773 ( .B1(n14735), .B2(n15761), .C1(n14783), .C2(n15519), .A(
        n2393), .ZN(n2390) );
  OAI22_X1 U774 ( .A1(n14667), .A2(n14845), .B1(n2287), .B2(n2288), .ZN(N975)
         );
  AOI221_X1 U775 ( .B1(n2297), .B2(n2298), .C1(n2299), .C2(n2300), .A(n14619), 
        .ZN(n2287) );
  AOI221_X1 U776 ( .B1(n2289), .B2(n2290), .C1(n2291), .C2(n2292), .A(n15293), 
        .ZN(n2288) );
  AOI221_X1 U777 ( .B1(n14735), .B2(n15760), .C1(n14783), .C2(n15518), .A(
        n2302), .ZN(n2299) );
  OAI22_X1 U778 ( .A1(n14697), .A2(n14845), .B1(n2062), .B2(n2068), .ZN(N985)
         );
  AOI221_X1 U779 ( .B1(n2085), .B2(n2086), .C1(n2087), .C2(n2088), .A(n14619), 
        .ZN(n2062) );
  AOI221_X1 U780 ( .B1(n2070), .B2(n2071), .C1(n2072), .C2(n2074), .A(n15293), 
        .ZN(n2068) );
  AOI221_X1 U781 ( .B1(n14734), .B2(n15758), .C1(n14783), .C2(n15516), .A(
        n2090), .ZN(n2087) );
  OAI22_X1 U782 ( .A1(n14700), .A2(n14845), .B1(n1938), .B2(n1942), .ZN(N986)
         );
  AOI221_X1 U783 ( .B1(n1975), .B2(n1976), .C1(n1978), .C2(n1982), .A(n14619), 
        .ZN(n1938) );
  AOI221_X1 U784 ( .B1(n1945), .B2(n1952), .C1(n1953), .C2(n1954), .A(n15293), 
        .ZN(n1942) );
  AOI221_X1 U785 ( .B1(n14734), .B2(n15757), .C1(n14783), .C2(n15515), .A(
        n2055), .ZN(n1978) );
  OAI22_X1 U786 ( .A1(n14703), .A2(n14845), .B1(n1861), .B2(n1862), .ZN(N987)
         );
  AOI221_X1 U787 ( .B1(n1877), .B2(n1881), .C1(n1883), .C2(n1884), .A(n14619), 
        .ZN(n1861) );
  AOI221_X1 U788 ( .B1(n1864), .B2(n1865), .C1(n1866), .C2(n1867), .A(n15293), 
        .ZN(n1862) );
  AOI221_X1 U789 ( .B1(n14733), .B2(n15756), .C1(n14783), .C2(n15514), .A(
        n1888), .ZN(n1883) );
  NAND2_X1 U790 ( .A1(n15302), .A2(n15301), .ZN(n1663) );
  BUF_X1 U791 ( .A(n1658), .Z(n14779) );
  BUF_X1 U792 ( .A(n1658), .Z(n14780) );
  INV_X1 U793 ( .A(n14828), .ZN(n14843) );
  INV_X1 U794 ( .A(n14716), .ZN(n14728) );
  NOR2_X1 U795 ( .A1(n2322), .A2(n15270), .ZN(n2180) );
  INV_X1 U796 ( .A(n2322), .ZN(n15293) );
  INV_X1 U797 ( .A(n2154), .ZN(n15289) );
  AND2_X1 U798 ( .A1(n2148), .A2(n14845), .ZN(n2564) );
  BUF_X1 U799 ( .A(n15294), .Z(n14618) );
  BUF_X1 U800 ( .A(n15294), .Z(n14619) );
  AOI21_X1 U801 ( .B1(n14842), .B2(n15730), .A(n15269), .ZN(n2550) );
  BUF_X1 U802 ( .A(n15267), .Z(n15274) );
  BUF_X1 U803 ( .A(n15266), .Z(n15272) );
  BUF_X1 U804 ( .A(n15266), .Z(n15273) );
  BUF_X1 U805 ( .A(n15267), .Z(n15275) );
  BUF_X1 U806 ( .A(n15266), .Z(n15271) );
  BUF_X1 U807 ( .A(n15267), .Z(n15276) );
  BUF_X1 U808 ( .A(n15268), .Z(n15277) );
  BUF_X1 U809 ( .A(n15268), .Z(n15278) );
  INV_X1 U810 ( .A(n14758), .ZN(n14774) );
  INV_X1 U811 ( .A(n14794), .ZN(n14810) );
  INV_X1 U812 ( .A(n1639), .ZN(n14827) );
  NOR3_X1 U813 ( .A1(n15282), .A2(n15283), .A3(n15284), .ZN(n3032) );
  NAND2_X1 U814 ( .A1(n2874), .A2(n2875), .ZN(N1008) );
  NOR4_X1 U815 ( .A1(n2884), .A2(n2885), .A3(n2886), .A4(n2887), .ZN(n2874) );
  NOR4_X1 U816 ( .A1(n2876), .A2(n2877), .A3(n2878), .A4(n2879), .ZN(n2875) );
  OAI221_X1 U817 ( .B1(n16183), .B2(n14860), .C1(n16114), .C2(n14857), .A(
        n2891), .ZN(n2884) );
  NAND2_X1 U818 ( .A1(n2856), .A2(n2857), .ZN(N1009) );
  NOR4_X1 U819 ( .A1(n2866), .A2(n2867), .A3(n2868), .A4(n2869), .ZN(n2856) );
  NOR4_X1 U820 ( .A1(n2858), .A2(n2859), .A3(n2860), .A4(n2861), .ZN(n2857) );
  OAI221_X1 U821 ( .B1(n16265), .B2(n14860), .C1(n16036), .C2(n14857), .A(
        n2873), .ZN(n2866) );
  NAND2_X1 U822 ( .A1(n2838), .A2(n2839), .ZN(N1010) );
  NOR4_X1 U823 ( .A1(n2848), .A2(n2849), .A3(n2850), .A4(n2851), .ZN(n2838) );
  NOR4_X1 U824 ( .A1(n2840), .A2(n2841), .A3(n2842), .A4(n2843), .ZN(n2839) );
  OAI221_X1 U825 ( .B1(n16172), .B2(n14860), .C1(n16113), .C2(n14857), .A(
        n2855), .ZN(n2848) );
  NAND2_X1 U826 ( .A1(n2820), .A2(n2821), .ZN(N1011) );
  NOR4_X1 U827 ( .A1(n2830), .A2(n2831), .A3(n2832), .A4(n2833), .ZN(n2820) );
  NOR4_X1 U828 ( .A1(n2822), .A2(n2823), .A3(n2824), .A4(n2825), .ZN(n2821) );
  OAI221_X1 U829 ( .B1(n16203), .B2(n14860), .C1(n16112), .C2(n14857), .A(
        n2837), .ZN(n2830) );
  NAND2_X1 U830 ( .A1(n2802), .A2(n2803), .ZN(N1012) );
  NOR4_X1 U831 ( .A1(n2812), .A2(n2813), .A3(n2814), .A4(n2815), .ZN(n2802) );
  NOR4_X1 U832 ( .A1(n2804), .A2(n2805), .A3(n2806), .A4(n2807), .ZN(n2803) );
  OAI221_X1 U833 ( .B1(n16182), .B2(n14861), .C1(n16111), .C2(n14858), .A(
        n2819), .ZN(n2812) );
  NAND2_X1 U834 ( .A1(n2784), .A2(n2785), .ZN(N1013) );
  NOR4_X1 U835 ( .A1(n2794), .A2(n2795), .A3(n2796), .A4(n2797), .ZN(n2784) );
  NOR4_X1 U836 ( .A1(n2786), .A2(n2787), .A3(n2788), .A4(n2789), .ZN(n2785) );
  OAI221_X1 U837 ( .B1(n16192), .B2(n14861), .C1(n15957), .C2(n14858), .A(
        n2801), .ZN(n2794) );
  NAND2_X1 U838 ( .A1(n2766), .A2(n2767), .ZN(N1014) );
  NOR4_X1 U839 ( .A1(n2776), .A2(n2777), .A3(n2778), .A4(n2779), .ZN(n2766) );
  NOR4_X1 U840 ( .A1(n2768), .A2(n2769), .A3(n2770), .A4(n2771), .ZN(n2767) );
  OAI221_X1 U841 ( .B1(n16191), .B2(n14861), .C1(n15956), .C2(n14858), .A(
        n2783), .ZN(n2776) );
  NAND2_X1 U842 ( .A1(n2748), .A2(n2749), .ZN(N1015) );
  NOR4_X1 U843 ( .A1(n2758), .A2(n2759), .A3(n2760), .A4(n2761), .ZN(n2748) );
  NOR4_X1 U844 ( .A1(n2750), .A2(n2751), .A3(n2752), .A4(n2753), .ZN(n2749) );
  OAI221_X1 U845 ( .B1(n16202), .B2(n14861), .C1(n16110), .C2(n14858), .A(
        n2765), .ZN(n2758) );
  NAND2_X1 U846 ( .A1(n2730), .A2(n2731), .ZN(N1016) );
  NOR4_X1 U847 ( .A1(n2740), .A2(n2741), .A3(n2742), .A4(n2743), .ZN(n2730) );
  NOR4_X1 U848 ( .A1(n2732), .A2(n2733), .A3(n2734), .A4(n2735), .ZN(n2731) );
  OAI221_X1 U849 ( .B1(n16264), .B2(n14861), .C1(n16035), .C2(n14858), .A(
        n2747), .ZN(n2740) );
  NAND2_X1 U850 ( .A1(n2712), .A2(n2713), .ZN(N1017) );
  NOR4_X1 U851 ( .A1(n2722), .A2(n2723), .A3(n2724), .A4(n2725), .ZN(n2712) );
  NOR4_X1 U852 ( .A1(n2714), .A2(n2715), .A3(n2716), .A4(n2717), .ZN(n2713) );
  OAI221_X1 U853 ( .B1(n16201), .B2(n14861), .C1(n16109), .C2(n14858), .A(
        n2729), .ZN(n2722) );
  NAND2_X1 U854 ( .A1(n2694), .A2(n2695), .ZN(N1018) );
  NOR4_X1 U855 ( .A1(n2704), .A2(n2705), .A3(n2706), .A4(n2707), .ZN(n2694) );
  NOR4_X1 U856 ( .A1(n2696), .A2(n2697), .A3(n2698), .A4(n2699), .ZN(n2695) );
  OAI221_X1 U857 ( .B1(n16181), .B2(n14861), .C1(n16108), .C2(n14858), .A(
        n2711), .ZN(n2704) );
  NAND2_X1 U858 ( .A1(n2676), .A2(n2677), .ZN(N1019) );
  NOR4_X1 U859 ( .A1(n2686), .A2(n2687), .A3(n2688), .A4(n2689), .ZN(n2676) );
  NOR4_X1 U860 ( .A1(n2678), .A2(n2679), .A3(n2680), .A4(n2681), .ZN(n2677) );
  OAI221_X1 U861 ( .B1(n16180), .B2(n14861), .C1(n16107), .C2(n14858), .A(
        n2693), .ZN(n2686) );
  NAND2_X1 U862 ( .A1(n2658), .A2(n2659), .ZN(N1020) );
  NOR4_X1 U863 ( .A1(n2668), .A2(n2669), .A3(n2670), .A4(n2671), .ZN(n2658) );
  NOR4_X1 U864 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659) );
  OAI221_X1 U865 ( .B1(n16179), .B2(n14861), .C1(n16106), .C2(n14858), .A(
        n2675), .ZN(n2668) );
  NAND2_X1 U866 ( .A1(n2640), .A2(n2641), .ZN(N1021) );
  NOR4_X1 U867 ( .A1(n2650), .A2(n2651), .A3(n2652), .A4(n2653), .ZN(n2640) );
  NOR4_X1 U868 ( .A1(n2642), .A2(n2643), .A3(n2644), .A4(n2645), .ZN(n2641) );
  OAI221_X1 U869 ( .B1(n16200), .B2(n14861), .C1(n16105), .C2(n14858), .A(
        n2657), .ZN(n2650) );
  NAND2_X1 U870 ( .A1(n2622), .A2(n2623), .ZN(N1022) );
  NOR4_X1 U871 ( .A1(n2632), .A2(n2633), .A3(n2634), .A4(n2635), .ZN(n2622) );
  NOR4_X1 U872 ( .A1(n2624), .A2(n2625), .A3(n2626), .A4(n2627), .ZN(n2623) );
  OAI221_X1 U873 ( .B1(n16293), .B2(n14861), .C1(n16039), .C2(n14858), .A(
        n2639), .ZN(n2632) );
  NAND2_X1 U874 ( .A1(n2604), .A2(n2605), .ZN(N1023) );
  NOR4_X1 U875 ( .A1(n2614), .A2(n2615), .A3(n2616), .A4(n2617), .ZN(n2604) );
  NOR4_X1 U876 ( .A1(n2606), .A2(n2607), .A3(n2608), .A4(n2609), .ZN(n2605) );
  OAI221_X1 U877 ( .B1(n16292), .B2(n14861), .C1(n16013), .C2(n14858), .A(
        n2621), .ZN(n2614) );
  NAND2_X1 U878 ( .A1(n1413), .A2(n1414), .ZN(N993) );
  NOR4_X1 U879 ( .A1(n1426), .A2(n1427), .A3(n1428), .A4(n1429), .ZN(n1413) );
  NOR4_X1 U880 ( .A1(n1415), .A2(n1416), .A3(n1417), .A4(n1418), .ZN(n1414) );
  OAI221_X1 U881 ( .B1(n16205), .B2(n14862), .C1(n16119), .C2(n14859), .A(
        n1435), .ZN(n1426) );
  NAND2_X1 U882 ( .A1(n1338), .A2(n1339), .ZN(N994) );
  NOR4_X1 U883 ( .A1(n1392), .A2(n1393), .A3(n1395), .A4(n1397), .ZN(n1338) );
  NOR4_X1 U884 ( .A1(n1340), .A2(n1341), .A3(n1342), .A4(n1344), .ZN(n1339) );
  OAI221_X1 U885 ( .B1(n16305), .B2(n14862), .C1(n16045), .C2(n14859), .A(
        n1412), .ZN(n1392) );
  NAND2_X1 U886 ( .A1(n1308), .A2(n1309), .ZN(N995) );
  NOR4_X1 U887 ( .A1(n1321), .A2(n1322), .A3(n1324), .A4(n1329), .ZN(n1308) );
  NOR4_X1 U888 ( .A1(n1310), .A2(n1311), .A3(n1312), .A4(n1313), .ZN(n1309) );
  OAI221_X1 U889 ( .B1(n16187), .B2(n14862), .C1(n16118), .C2(n14859), .A(
        n1336), .ZN(n1321) );
  NAND2_X1 U890 ( .A1(n1287), .A2(n1288), .ZN(N996) );
  NOR4_X1 U891 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1287) );
  NOR4_X1 U892 ( .A1(n1289), .A2(n1290), .A3(n1291), .A4(n1292), .ZN(n1288) );
  OAI221_X1 U893 ( .B1(n16304), .B2(n14862), .C1(n16117), .C2(n14859), .A(
        n1307), .ZN(n1299) );
  NAND2_X1 U894 ( .A1(n1258), .A2(n1260), .ZN(N997) );
  NOR4_X1 U895 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1258) );
  NOR4_X1 U896 ( .A1(n1265), .A2(n1268), .A3(n1269), .A4(n1272), .ZN(n1260) );
  OAI221_X1 U897 ( .B1(n16254), .B2(n14862), .C1(n16044), .C2(n14859), .A(
        n1286), .ZN(n1278) );
  NAND2_X1 U898 ( .A1(n1209), .A2(n1211), .ZN(N998) );
  NOR4_X1 U899 ( .A1(n1232), .A2(n1234), .A3(n1239), .A4(n1241), .ZN(n1209) );
  NOR4_X1 U900 ( .A1(n1212), .A2(n1213), .A3(n1222), .A4(n1224), .ZN(n1211) );
  OAI221_X1 U901 ( .B1(n16204), .B2(n14862), .C1(n16116), .C2(n14859), .A(
        n1257), .ZN(n1232) );
  NAND2_X1 U902 ( .A1(n1128), .A2(n1129), .ZN(N999) );
  NOR4_X1 U903 ( .A1(n1154), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1128) );
  NOR4_X1 U904 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
  OAI221_X1 U905 ( .B1(n16253), .B2(n14862), .C1(n16043), .C2(n14859), .A(
        n1201), .ZN(n1154) );
  NAND2_X1 U906 ( .A1(n2586), .A2(n2587), .ZN(N1024) );
  NOR4_X1 U907 ( .A1(n2596), .A2(n2597), .A3(n2598), .A4(n2599), .ZN(n2586) );
  NOR4_X1 U908 ( .A1(n2588), .A2(n2589), .A3(n2590), .A4(n2591), .ZN(n2587) );
  OAI221_X1 U909 ( .B1(n16291), .B2(n14862), .C1(n16012), .C2(n14859), .A(
        n2603), .ZN(n2596) );
  OAI221_X1 U910 ( .B1(n16015), .B2(n14932), .C1(n15566), .C2(n14929), .A(
        n2863), .ZN(n2860) );
  AOI22_X1 U911 ( .A1(n14926), .A2(n15488), .B1(n14924), .B2(n15416), .ZN(
        n2863) );
  OAI221_X1 U912 ( .B1(n16014), .B2(n14933), .C1(n15565), .C2(n14930), .A(
        n2737), .ZN(n2734) );
  AOI22_X1 U913 ( .A1(n14927), .A2(n15485), .B1(n14924), .B2(n15411), .ZN(
        n2737) );
  NAND2_X1 U914 ( .A1(n3038), .A2(n3029), .ZN(n1150) );
  NAND2_X1 U915 ( .A1(n3038), .A2(n3026), .ZN(n1161) );
  NAND2_X1 U916 ( .A1(n3036), .A2(n3029), .ZN(n1145) );
  NAND2_X1 U917 ( .A1(n3025), .A2(n3029), .ZN(n1134) );
  NAND2_X1 U918 ( .A1(n3025), .A2(n3028), .ZN(n1135) );
  NAND2_X1 U919 ( .A1(n3028), .A2(n3038), .ZN(n1144) );
  NAND2_X1 U920 ( .A1(n3027), .A2(n3038), .ZN(n1170) );
  NAND2_X1 U921 ( .A1(n3032), .A2(n3038), .ZN(n1160) );
  NAND2_X1 U922 ( .A1(n3033), .A2(n3038), .ZN(n1178) );
  NAND2_X1 U923 ( .A1(n3031), .A2(n3036), .ZN(n1168) );
  NAND2_X1 U924 ( .A1(n3033), .A2(n3036), .ZN(n1196) );
  NAND2_X1 U925 ( .A1(n3034), .A2(n3025), .ZN(n1139) );
  NAND2_X1 U926 ( .A1(n3033), .A2(n3025), .ZN(n1140) );
  NAND2_X1 U927 ( .A1(n3026), .A2(n3037), .ZN(n1149) );
  NAND2_X1 U928 ( .A1(n3034), .A2(n3037), .ZN(n1194) );
  OAI22_X1 U929 ( .A1(n15263), .A2(n14653), .B1(n15258), .B2(n16313), .ZN(
        n2125) );
  OAI22_X1 U930 ( .A1(n15263), .A2(n14656), .B1(n15258), .B2(n16312), .ZN(
        n2126) );
  OAI22_X1 U931 ( .A1(n15262), .A2(n14683), .B1(n15258), .B2(n16311), .ZN(
        n2135) );
  OAI22_X1 U932 ( .A1(n15264), .A2(n14641), .B1(n15257), .B2(n16306), .ZN(
        n2121) );
  OAI22_X1 U933 ( .A1(n15265), .A2(n14620), .B1(n15257), .B2(n16290), .ZN(
        n2114) );
  OAI22_X1 U934 ( .A1(n15264), .A2(n14635), .B1(n15258), .B2(n16289), .ZN(
        n2119) );
  OAI22_X1 U935 ( .A1(n15263), .A2(n14674), .B1(n15258), .B2(n16288), .ZN(
        n2132) );
  OAI22_X1 U936 ( .A1(n15262), .A2(n14686), .B1(n15258), .B2(n16287), .ZN(
        n2136) );
  OAI22_X1 U937 ( .A1(n15262), .A2(n14692), .B1(n15258), .B2(n16286), .ZN(
        n2138) );
  OAI22_X1 U938 ( .A1(n15261), .A2(n14704), .B1(n15258), .B2(n16285), .ZN(
        n2142) );
  OAI22_X1 U939 ( .A1(n15261), .A2(n14710), .B1(n15257), .B2(n16284), .ZN(
        n2144) );
  OAI22_X1 U940 ( .A1(n15260), .A2(n14713), .B1(n15257), .B2(n16283), .ZN(
        n2145) );
  OAI22_X1 U941 ( .A1(n15259), .A2(n14671), .B1(n15257), .B2(n16263), .ZN(
        n3625) );
  OAI22_X1 U942 ( .A1(n15261), .A2(n14707), .B1(n15257), .B2(n16262), .ZN(
        n2143) );
  OAI22_X1 U943 ( .A1(n15259), .A2(n14632), .B1(n15257), .B2(n16252), .ZN(
        n3609) );
  OAI22_X1 U944 ( .A1(n15260), .A2(n14638), .B1(n15257), .B2(n16251), .ZN(
        n3388) );
  OAI22_X1 U945 ( .A1(n15259), .A2(n14647), .B1(n15257), .B2(n16250), .ZN(
        n3608) );
  OAI22_X1 U946 ( .A1(n15260), .A2(n14662), .B1(n15257), .B2(n16249), .ZN(
        n3387) );
  OAI22_X1 U947 ( .A1(n15260), .A2(n14668), .B1(n15257), .B2(n16248), .ZN(
        n3386) );
  OAI22_X1 U948 ( .A1(n15260), .A2(n14689), .B1(n15257), .B2(n16247), .ZN(
        n3385) );
  OAI22_X1 U949 ( .A1(n15264), .A2(n14626), .B1(n15257), .B2(n16227), .ZN(
        n2116) );
  OAI22_X1 U950 ( .A1(n15264), .A2(n14629), .B1(n15258), .B2(n16226), .ZN(
        n2117) );
  OAI22_X1 U951 ( .A1(n15264), .A2(n14650), .B1(n15257), .B2(n16225), .ZN(
        n2124) );
  OAI22_X1 U952 ( .A1(n15263), .A2(n14665), .B1(n15258), .B2(n16224), .ZN(
        n2129) );
  OAI22_X1 U953 ( .A1(n15263), .A2(n14677), .B1(n15258), .B2(n16223), .ZN(
        n2133) );
  OAI22_X1 U954 ( .A1(n15262), .A2(n14695), .B1(n15258), .B2(n16222), .ZN(
        n2139) );
  OAI22_X1 U955 ( .A1(n15261), .A2(n14698), .B1(n15258), .B2(n16221), .ZN(
        n2140) );
  OAI22_X1 U956 ( .A1(n15261), .A2(n14701), .B1(n15258), .B2(n16220), .ZN(
        n2141) );
  OAI22_X1 U957 ( .A1(n15265), .A2(n14623), .B1(n15258), .B2(n16207), .ZN(
        n2115) );
  OAI22_X1 U958 ( .A1(n15259), .A2(n14659), .B1(n15257), .B2(n16206), .ZN(
        n3626) );
  OAI22_X1 U959 ( .A1(n15262), .A2(n14680), .B1(n15258), .B2(n16199), .ZN(
        n2134) );
  OAI22_X1 U960 ( .A1(n14655), .A2(n1126), .B1(n14953), .B2(n15785), .ZN(n1357) );
  OAI22_X1 U961 ( .A1(n14658), .A2(n1126), .B1(n14952), .B2(n15784), .ZN(n1358) );
  OAI22_X1 U962 ( .A1(n14682), .A2(n1126), .B1(n14950), .B2(n15783), .ZN(n1366) );
  OAI22_X1 U963 ( .A1(n14685), .A2(n14947), .B1(n14950), .B2(n15782), .ZN(
        n1367) );
  OAI22_X1 U964 ( .A1(n14652), .A2(n1126), .B1(n14953), .B2(n15761), .ZN(n1356) );
  OAI22_X1 U965 ( .A1(n14667), .A2(n1126), .B1(n14952), .B2(n15760), .ZN(n1361) );
  OAI22_X1 U966 ( .A1(n14679), .A2(n1126), .B1(n14951), .B2(n15759), .ZN(n1365) );
  OAI22_X1 U967 ( .A1(n14697), .A2(n1126), .B1(n14949), .B2(n15758), .ZN(n1371) );
  OAI22_X1 U968 ( .A1(n14700), .A2(n14947), .B1(n14949), .B2(n15757), .ZN(
        n1372) );
  OAI22_X1 U969 ( .A1(n14703), .A2(n14947), .B1(n14949), .B2(n15756), .ZN(
        n1373) );
  OAI22_X1 U970 ( .A1(n14670), .A2(n1126), .B1(n14951), .B2(n15752), .ZN(n1362) );
  OAI22_X1 U971 ( .A1(n14691), .A2(n1126), .B1(n14950), .B2(n15751), .ZN(n1369) );
  OAI22_X1 U972 ( .A1(n14628), .A2(n1126), .B1(n14955), .B2(n15649), .ZN(n1348) );
  OAI22_X1 U973 ( .A1(n14631), .A2(n1126), .B1(n14955), .B2(n15648), .ZN(n1349) );
  OAI22_X1 U974 ( .A1(n14643), .A2(n1126), .B1(n14954), .B2(n15647), .ZN(n1353) );
  OAI22_X1 U975 ( .A1(n14673), .A2(n1126), .B1(n14951), .B2(n15607), .ZN(n1363) );
  OAI22_X1 U976 ( .A1(n14634), .A2(n1126), .B1(n14954), .B2(n15578), .ZN(n1350) );
  OAI22_X1 U977 ( .A1(n14640), .A2(n1126), .B1(n14954), .B2(n15577), .ZN(n1352) );
  OAI22_X1 U978 ( .A1(n14649), .A2(n1126), .B1(n14953), .B2(n15576), .ZN(n1355) );
  OAI22_X1 U979 ( .A1(n14664), .A2(n1126), .B1(n14952), .B2(n15575), .ZN(n1360) );
  OAI22_X1 U980 ( .A1(n14625), .A2(n14947), .B1(n14955), .B2(n15542), .ZN(
        n1347) );
  OAI22_X1 U981 ( .A1(n14661), .A2(n1126), .B1(n14952), .B2(n15541), .ZN(n1359) );
  OAI22_X1 U982 ( .A1(n14712), .A2(n1126), .B1(n14948), .B2(n15538), .ZN(n1376) );
  OAI22_X1 U983 ( .A1(n14715), .A2(n1126), .B1(n14948), .B2(n15537), .ZN(n1377) );
  AND2_X1 U984 ( .A1(n3036), .A2(n3026), .ZN(n1152) );
  AND2_X1 U985 ( .A1(n3025), .A2(n3026), .ZN(n1138) );
  AND2_X1 U986 ( .A1(n3034), .A2(n3038), .ZN(n1202) );
  AND2_X1 U987 ( .A1(n3028), .A2(n3036), .ZN(n1148) );
  AND2_X1 U988 ( .A1(n3034), .A2(n3036), .ZN(n1176) );
  AND2_X1 U989 ( .A1(n3027), .A2(n3036), .ZN(n1163) );
  AND2_X1 U990 ( .A1(n3027), .A2(n3025), .ZN(n1137) );
  AND2_X1 U991 ( .A1(n3031), .A2(n3025), .ZN(n1143) );
  AND2_X1 U992 ( .A1(n3032), .A2(n3025), .ZN(n1142) );
  AND2_X1 U993 ( .A1(n3028), .A2(n3037), .ZN(n1147) );
  AND2_X1 U994 ( .A1(n3029), .A2(n3037), .ZN(n1153) );
  AND2_X1 U995 ( .A1(n3027), .A2(n3037), .ZN(n1172) );
  AND2_X1 U996 ( .A1(n3031), .A2(n3037), .ZN(n1189) );
  AND2_X1 U997 ( .A1(n3032), .A2(n3037), .ZN(n1188) );
  AND2_X1 U998 ( .A1(n3033), .A2(n3037), .ZN(n1205) );
  NAND2_X1 U999 ( .A1(n3018), .A2(n3019), .ZN(N1000) );
  NOR4_X1 U1000 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n3018)
         );
  NOR4_X1 U1001 ( .A1(n3020), .A2(n3021), .A3(n3022), .A4(n3023), .ZN(n3019)
         );
  OAI221_X1 U1002 ( .B1(n16244), .B2(n14860), .C1(n16089), .C2(n14857), .A(
        n3047), .ZN(n3040) );
  NAND2_X1 U1003 ( .A1(n3000), .A2(n3001), .ZN(N1001) );
  NOR4_X1 U1004 ( .A1(n3010), .A2(n3011), .A3(n3012), .A4(n3013), .ZN(n3000)
         );
  NOR4_X1 U1005 ( .A1(n3002), .A2(n3003), .A3(n3004), .A4(n3005), .ZN(n3001)
         );
  OAI221_X1 U1006 ( .B1(n16294), .B2(n14860), .C1(n16088), .C2(n14857), .A(
        n3017), .ZN(n3010) );
  NAND2_X1 U1007 ( .A1(n2982), .A2(n2983), .ZN(N1002) );
  NOR4_X1 U1008 ( .A1(n2992), .A2(n2993), .A3(n2994), .A4(n2995), .ZN(n2982)
         );
  NOR4_X1 U1009 ( .A1(n2984), .A2(n2985), .A3(n2986), .A4(n2987), .ZN(n2983)
         );
  OAI221_X1 U1010 ( .B1(n16186), .B2(n14860), .C1(n16042), .C2(n14857), .A(
        n2999), .ZN(n2992) );
  NAND2_X1 U1011 ( .A1(n2964), .A2(n2965), .ZN(N1003) );
  NOR4_X1 U1012 ( .A1(n2974), .A2(n2975), .A3(n2976), .A4(n2977), .ZN(n2964)
         );
  NOR4_X1 U1013 ( .A1(n2966), .A2(n2967), .A3(n2968), .A4(n2969), .ZN(n2965)
         );
  OAI221_X1 U1014 ( .B1(n16185), .B2(n14860), .C1(n16115), .C2(n14857), .A(
        n2981), .ZN(n2974) );
  NAND2_X1 U1015 ( .A1(n2946), .A2(n2947), .ZN(N1004) );
  NOR4_X1 U1016 ( .A1(n2956), .A2(n2957), .A3(n2958), .A4(n2959), .ZN(n2946)
         );
  NOR4_X1 U1017 ( .A1(n2948), .A2(n2949), .A3(n2950), .A4(n2951), .ZN(n2947)
         );
  OAI221_X1 U1018 ( .B1(n16194), .B2(n14860), .C1(n15959), .C2(n14857), .A(
        n2963), .ZN(n2956) );
  NAND2_X1 U1019 ( .A1(n2928), .A2(n2929), .ZN(N1005) );
  NOR4_X1 U1020 ( .A1(n2938), .A2(n2939), .A3(n2940), .A4(n2941), .ZN(n2928)
         );
  NOR4_X1 U1021 ( .A1(n2930), .A2(n2931), .A3(n2932), .A4(n2933), .ZN(n2929)
         );
  OAI221_X1 U1022 ( .B1(n16193), .B2(n14860), .C1(n15958), .C2(n14857), .A(
        n2945), .ZN(n2938) );
  NAND2_X1 U1023 ( .A1(n2910), .A2(n2911), .ZN(N1006) );
  NOR4_X1 U1024 ( .A1(n2920), .A2(n2921), .A3(n2922), .A4(n2923), .ZN(n2910)
         );
  NOR4_X1 U1025 ( .A1(n2912), .A2(n2913), .A3(n2914), .A4(n2915), .ZN(n2911)
         );
  OAI221_X1 U1026 ( .B1(n16184), .B2(n14860), .C1(n16041), .C2(n14857), .A(
        n2927), .ZN(n2920) );
  NAND2_X1 U1027 ( .A1(n2892), .A2(n2893), .ZN(N1007) );
  NOR4_X1 U1028 ( .A1(n2902), .A2(n2903), .A3(n2904), .A4(n2905), .ZN(n2892)
         );
  NOR4_X1 U1029 ( .A1(n2894), .A2(n2895), .A3(n2896), .A4(n2897), .ZN(n2893)
         );
  OAI221_X1 U1030 ( .B1(n16296), .B2(n14860), .C1(n16040), .C2(n14857), .A(
        n2909), .ZN(n2902) );
  OAI22_X1 U1031 ( .A1(n15110), .A2(n16305), .B1(n15108), .B2(n14623), .ZN(
        n3429) );
  OAI22_X1 U1032 ( .A1(n15116), .A2(n16304), .B1(n14630), .B2(n15108), .ZN(
        n1701) );
  OAI22_X1 U1033 ( .A1(n15115), .A2(n16294), .B1(n14645), .B2(n15109), .ZN(
        n1706) );
  OAI22_X1 U1034 ( .A1(n15112), .A2(n16293), .B1(n14708), .B2(n15108), .ZN(
        n3419) );
  OAI22_X1 U1035 ( .A1(n15247), .A2(n16269), .B1(n15251), .B2(n14707), .ZN(
        n2079) );
  OAI22_X1 U1036 ( .A1(n15138), .A2(n16267), .B1(n14641), .B2(n15135), .ZN(
        n3585) );
  OAI22_X1 U1037 ( .A1(n15139), .A2(n16266), .B1(n14644), .B2(n15135), .ZN(
        n3584) );
  OAI22_X1 U1038 ( .A1(n15110), .A2(n16254), .B1(n14633), .B2(n15108), .ZN(
        n3428) );
  OAI22_X1 U1039 ( .A1(n15111), .A2(n16253), .B1(n14639), .B2(n15108), .ZN(
        n3426) );
  OAI22_X1 U1040 ( .A1(n15247), .A2(n16235), .B1(n15251), .B2(n14710), .ZN(
        n2080) );
  OAI22_X1 U1041 ( .A1(n15247), .A2(n16234), .B1(n15250), .B2(n14713), .ZN(
        n2081) );
  OAI22_X1 U1042 ( .A1(n15247), .A2(n16229), .B1(n15255), .B2(n14623), .ZN(
        n2051) );
  OAI22_X1 U1043 ( .A1(n15137), .A2(n16190), .B1(n14665), .B2(n15135), .ZN(
        n3618) );
  OAI22_X1 U1044 ( .A1(n15116), .A2(n16187), .B1(n14627), .B2(n15108), .ZN(
        n1700) );
  OAI22_X1 U1045 ( .A1(n15115), .A2(n16186), .B1(n14648), .B2(n15108), .ZN(
        n1707) );
  OAI22_X1 U1046 ( .A1(n15115), .A2(n16185), .B1(n14651), .B2(n15109), .ZN(
        n1708) );
  OAI22_X1 U1047 ( .A1(n15114), .A2(n16183), .B1(n14666), .B2(n15109), .ZN(
        n1713) );
  OAI22_X1 U1048 ( .A1(n15114), .A2(n16182), .B1(n14678), .B2(n15109), .ZN(
        n1717) );
  OAI22_X1 U1049 ( .A1(n15113), .A2(n16181), .B1(n14696), .B2(n15109), .ZN(
        n1723) );
  OAI22_X1 U1050 ( .A1(n15113), .A2(n16180), .B1(n14699), .B2(n15109), .ZN(
        n1724) );
  OAI22_X1 U1051 ( .A1(n15113), .A2(n16179), .B1(n14702), .B2(n15109), .ZN(
        n1725) );
  OAI22_X1 U1052 ( .A1(n15121), .A2(n16178), .B1(n14645), .B2(n15117), .ZN(
        n3463) );
  OAI22_X1 U1053 ( .A1(n15111), .A2(n16172), .B1(n14672), .B2(n15108), .ZN(
        n3424) );
  OAI22_X1 U1054 ( .A1(n15054), .A2(n16169), .B1(n14641), .B2(n15050), .ZN(
        n3507) );
  OAI22_X1 U1055 ( .A1(n15055), .A2(n16168), .B1(n14673), .B2(n15050), .ZN(
        n3501) );
  OAI22_X1 U1056 ( .A1(n15123), .A2(n16167), .B1(n14671), .B2(n15118), .ZN(
        n1331) );
  OAI22_X1 U1057 ( .A1(n15235), .A2(n16153), .B1(n1081), .B2(n14641), .ZN(
        n3598) );
  OAI22_X1 U1058 ( .A1(n15235), .A2(n16152), .B1(n14644), .B2(n15233), .ZN(
        n3597) );
  OAI22_X1 U1059 ( .A1(n15236), .A2(n16104), .B1(n1081), .B2(n14647), .ZN(
        n3596) );
  OAI22_X1 U1060 ( .A1(n15246), .A2(n16103), .B1(n15255), .B2(n14632), .ZN(
        n2054) );
  OAI22_X1 U1061 ( .A1(n15246), .A2(n16102), .B1(n15254), .B2(n14638), .ZN(
        n2056) );
  OAI22_X1 U1062 ( .A1(n15247), .A2(n16101), .B1(n15253), .B2(n14671), .ZN(
        n2067) );
  OAI22_X1 U1063 ( .A1(n15235), .A2(n16087), .B1(n1081), .B2(n14629), .ZN(
        n3599) );
  OAI22_X1 U1064 ( .A1(n15132), .A2(n16048), .B1(n14666), .B2(n15127), .ZN(
        n1681) );
  OAI22_X1 U1065 ( .A1(n15131), .A2(n16047), .B1(n14678), .B2(n15127), .ZN(
        n1685) );
  OAI22_X1 U1066 ( .A1(n15130), .A2(n16046), .B1(n14696), .B2(n15127), .ZN(
        n1691) );
  OAI22_X1 U1067 ( .A1(n15151), .A2(n16009), .B1(n14642), .B2(n15145), .ZN(
        n1641) );
  OAI22_X1 U1068 ( .A1(n15151), .A2(n16008), .B1(n14645), .B2(n15144), .ZN(
        n1642) );
  OAI22_X1 U1069 ( .A1(n15134), .A2(n15960), .B1(n15127), .B2(n14623), .ZN(
        n1667) );
  OAI22_X1 U1070 ( .A1(n15128), .A2(n15950), .B1(n14711), .B2(n15126), .ZN(
        n3612) );
  OAI22_X1 U1071 ( .A1(n15128), .A2(n15949), .B1(n14713), .B2(n15126), .ZN(
        n3611) );
  OAI22_X1 U1072 ( .A1(n15028), .A2(n15948), .B1(n14621), .B2(n15020), .ZN(
        n1890) );
  OAI22_X1 U1073 ( .A1(n15027), .A2(n15946), .B1(n14636), .B2(n15020), .ZN(
        n1895) );
  OAI22_X1 U1074 ( .A1(n15024), .A2(n15942), .B1(n14672), .B2(n15021), .ZN(
        n1907) );
  OAI22_X1 U1075 ( .A1(n15024), .A2(n15941), .B1(n14675), .B2(n15021), .ZN(
        n1908) );
  OAI22_X1 U1076 ( .A1(n15023), .A2(n15940), .B1(n14687), .B2(n15021), .ZN(
        n1912) );
  OAI22_X1 U1077 ( .A1(n15023), .A2(n15939), .B1(n14693), .B2(n15020), .ZN(
        n1914) );
  OAI22_X1 U1078 ( .A1(n15022), .A2(n15938), .B1(n14705), .B2(n15021), .ZN(
        n1918) );
  OAI22_X1 U1079 ( .A1(n15022), .A2(n15937), .B1(n14708), .B2(n15020), .ZN(
        n1919) );
  OAI22_X1 U1080 ( .A1(n15046), .A2(n15916), .B1(n14654), .B2(n15040), .ZN(
        n2029) );
  OAI22_X1 U1081 ( .A1(n15044), .A2(n15914), .B1(n14680), .B2(n1110), .ZN(
        n2038) );
  OAI22_X1 U1082 ( .A1(n15043), .A2(n15892), .B1(n14708), .B2(n1110), .ZN(
        n2047) );
  OAI22_X1 U1083 ( .A1(n15037), .A2(n15885), .B1(n14627), .B2(n1112), .ZN(
        n1988) );
  OAI22_X1 U1084 ( .A1(n15037), .A2(n15884), .B1(n14630), .B2(n1112), .ZN(
        n1989) );
  OAI22_X1 U1085 ( .A1(n15036), .A2(n15882), .B1(n14644), .B2(n1112), .ZN(
        n1994) );
  OAI22_X1 U1086 ( .A1(n15036), .A2(n15881), .B1(n14651), .B2(n15029), .ZN(
        n1996) );
  OAI22_X1 U1087 ( .A1(n15035), .A2(n15880), .B1(n14666), .B2(n1112), .ZN(
        n2001) );
  OAI22_X1 U1088 ( .A1(n15034), .A2(n15877), .B1(n14678), .B2(n1112), .ZN(
        n2005) );
  OAI22_X1 U1089 ( .A1(n15033), .A2(n15875), .B1(n14696), .B2(n1112), .ZN(
        n2011) );
  OAI22_X1 U1090 ( .A1(n15034), .A2(n15874), .B1(n14699), .B2(n1112), .ZN(
        n2012) );
  OAI22_X1 U1091 ( .A1(n15033), .A2(n15873), .B1(n14702), .B2(n1112), .ZN(
        n2013) );
  OAI22_X1 U1092 ( .A1(n15036), .A2(n15847), .B1(n14648), .B2(n15029), .ZN(
        n1995) );
  OAI22_X1 U1093 ( .A1(n15197), .A2(n15845), .B1(n14648), .B2(n15200), .ZN(
        n1195) );
  OAI22_X1 U1094 ( .A1(n15169), .A2(n15830), .B1(n14643), .B2(n15164), .ZN(
        n1225) );
  OAI22_X1 U1095 ( .A1(n15095), .A2(n15821), .B1(n14667), .B2(n1095), .ZN(
        n1169) );
  OAI22_X1 U1096 ( .A1(n15095), .A2(n15820), .B1(n14679), .B2(n1095), .ZN(
        n1173) );
  OAI22_X1 U1097 ( .A1(n15095), .A2(n15819), .B1(n14697), .B2(n1095), .ZN(
        n1179) );
  OAI22_X1 U1098 ( .A1(n15073), .A2(n15795), .B1(n14664), .B2(n1097), .ZN(
        n3546) );
  OAI22_X1 U1099 ( .A1(n15179), .A2(n15697), .B1(n15174), .B2(n14713), .ZN(
        n1985) );
  OAI22_X1 U1100 ( .A1(n14966), .A2(n15684), .B1(n14620), .B2(n1125), .ZN(
        n1474) );
  OAI22_X1 U1101 ( .A1(n14966), .A2(n15683), .B1(n14628), .B2(n14958), .ZN(
        n1476) );
  OAI22_X1 U1102 ( .A1(n14962), .A2(n15681), .B1(n14674), .B2(n1125), .ZN(
        n1492) );
  OAI22_X1 U1103 ( .A1(n14960), .A2(n15679), .B1(n14692), .B2(n1125), .ZN(
        n1498) );
  OAI22_X1 U1104 ( .A1(n14959), .A2(n15677), .B1(n14709), .B2(n1125), .ZN(
        n1503) );
  OAI22_X1 U1105 ( .A1(n15198), .A2(n15668), .B1(n15206), .B2(n14624), .ZN(
        n1187) );
  OAI22_X1 U1106 ( .A1(n14986), .A2(n15651), .B1(n14647), .B2(n1123), .ZN(
        n1547) );
  OAI22_X1 U1107 ( .A1(n14984), .A2(n15586), .B1(n14669), .B2(n1123), .ZN(
        n1554) );
  OAI22_X1 U1108 ( .A1(n14982), .A2(n15584), .B1(n14690), .B2(n1123), .ZN(
        n1561) );
  OAI22_X1 U1109 ( .A1(n14987), .A2(n15583), .B1(n14630), .B2(n14979), .ZN(
        n1541) );
  OAI22_X1 U1110 ( .A1(n14966), .A2(n15531), .B1(n14625), .B2(n1125), .ZN(
        n1475) );
  OAI22_X1 U1111 ( .A1(n14964), .A2(n15519), .B1(n14652), .B2(n1125), .ZN(
        n1484) );
  OAI22_X1 U1112 ( .A1(n14963), .A2(n15518), .B1(n14667), .B2(n1125), .ZN(
        n1489) );
  OAI22_X1 U1113 ( .A1(n14962), .A2(n15517), .B1(n14679), .B2(n1125), .ZN(
        n1493) );
  OAI22_X1 U1114 ( .A1(n14960), .A2(n15516), .B1(n14697), .B2(n14958), .ZN(
        n1499) );
  OAI22_X1 U1115 ( .A1(n14960), .A2(n15515), .B1(n14700), .B2(n1125), .ZN(
        n1500) );
  OAI22_X1 U1116 ( .A1(n14964), .A2(n15505), .B1(n14648), .B2(n1125), .ZN(
        n1483) );
  OAI22_X1 U1117 ( .A1(n14962), .A2(n15434), .B1(n14670), .B2(n1125), .ZN(
        n1490) );
  OAI22_X1 U1118 ( .A1(n14961), .A2(n15433), .B1(n14691), .B2(n1125), .ZN(
        n1497) );
  OAI22_X1 U1119 ( .A1(n14966), .A2(n15426), .B1(n14631), .B2(n1125), .ZN(
        n1477) );
  OAI22_X1 U1120 ( .A1(n15115), .A2(n16244), .B1(n14642), .B2(n15109), .ZN(
        n1705) );
  OAI22_X1 U1121 ( .A1(n15247), .A2(n16228), .B1(n15255), .B2(n14629), .ZN(
        n2053) );
  OAI22_X1 U1122 ( .A1(n15112), .A2(n16201), .B1(n14693), .B2(n15108), .ZN(
        n3421) );
  OAI22_X1 U1123 ( .A1(n15112), .A2(n16200), .B1(n14705), .B2(n15108), .ZN(
        n3420) );
  OAI22_X1 U1124 ( .A1(n15137), .A2(n16189), .B1(n14678), .B2(n15135), .ZN(
        n3617) );
  OAI22_X1 U1125 ( .A1(n15137), .A2(n16188), .B1(n14695), .B2(n15135), .ZN(
        n3616) );
  OAI22_X1 U1126 ( .A1(n15122), .A2(n16174), .B1(n14709), .B2(n15118), .ZN(
        n1343) );
  OAI22_X1 U1127 ( .A1(n15236), .A2(n16151), .B1(n1081), .B2(n14659), .ZN(
        n3595) );
  OAI22_X1 U1128 ( .A1(n15026), .A2(n16066), .B1(n14654), .B2(n15020), .ZN(
        n1901) );
  OAI22_X1 U1129 ( .A1(n15025), .A2(n16065), .B1(n14657), .B2(n15021), .ZN(
        n1902) );
  OAI22_X1 U1130 ( .A1(n15024), .A2(n16063), .B1(n14681), .B2(n15021), .ZN(
        n1910) );
  OAI22_X1 U1131 ( .A1(n15024), .A2(n16062), .B1(n14684), .B2(n15021), .ZN(
        n1911) );
  OAI22_X1 U1132 ( .A1(n15025), .A2(n15943), .B1(n14663), .B2(n15021), .ZN(
        n1904) );
  OAI22_X1 U1133 ( .A1(n15046), .A2(n15915), .B1(n14657), .B2(n1110), .ZN(
        n2030) );
  OAI22_X1 U1134 ( .A1(n15044), .A2(n15913), .B1(n14684), .B2(n1110), .ZN(
        n2039) );
  OAI22_X1 U1135 ( .A1(n15046), .A2(n15899), .B1(n14660), .B2(n1110), .ZN(
        n2031) );
  OAI22_X1 U1136 ( .A1(n15180), .A2(n15860), .B1(n14660), .B2(n15174), .ZN(
        n1967) );
  OAI22_X1 U1137 ( .A1(n15094), .A2(n15853), .B1(n14680), .B2(n1095), .ZN(
        n1174) );
  OAI22_X1 U1138 ( .A1(n15177), .A2(n15698), .B1(n15174), .B2(n14710), .ZN(
        n1984) );
  OAI22_X1 U1139 ( .A1(n14965), .A2(n15682), .B1(n14635), .B2(n1125), .ZN(
        n1479) );
  OAI22_X1 U1140 ( .A1(n14959), .A2(n15678), .B1(n14704), .B2(n1125), .ZN(
        n1502) );
  OAI22_X1 U1141 ( .A1(n14960), .A2(n15514), .B1(n14703), .B2(n1125), .ZN(
        n1501) );
  OAI22_X1 U1142 ( .A1(n14963), .A2(n15497), .B1(n14715), .B2(n1125), .ZN(
        n1505) );
  OAI22_X1 U1143 ( .A1(n15111), .A2(n16296), .B1(n14663), .B2(n15108), .ZN(
        n3425) );
  OAI22_X1 U1144 ( .A1(n15143), .A2(n16257), .B1(n14647), .B2(n15135), .ZN(
        n1419) );
  OAI22_X1 U1145 ( .A1(n15124), .A2(n16177), .B1(n14661), .B2(n15118), .ZN(
        n1327) );
  OAI22_X1 U1146 ( .A1(n15123), .A2(n16176), .B1(n14670), .B2(n15118), .ZN(
        n1330) );
  OAI22_X1 U1147 ( .A1(n15123), .A2(n16175), .B1(n14691), .B2(n15118), .ZN(
        n1337) );
  OAI22_X1 U1148 ( .A1(n15057), .A2(n16171), .B1(n15050), .B2(n14623), .ZN(
        n3511) );
  OAI22_X1 U1149 ( .A1(n15246), .A2(n16149), .B1(n14644), .B2(n15248), .ZN(
        n2058) );
  OAI22_X1 U1150 ( .A1(n15133), .A2(n16095), .B1(n14630), .B2(n15126), .ZN(
        n1669) );
  OAI22_X1 U1151 ( .A1(n15133), .A2(n16038), .B1(n14648), .B2(n15127), .ZN(
        n1675) );
  OAI22_X1 U1152 ( .A1(n15132), .A2(n16037), .B1(n14660), .B2(n15127), .ZN(
        n1679) );
  OAI22_X1 U1153 ( .A1(n15027), .A2(n16023), .B1(n14627), .B2(n15020), .ZN(
        n1892) );
  OAI22_X1 U1154 ( .A1(n15026), .A2(n16021), .B1(n14651), .B2(n15020), .ZN(
        n1900) );
  OAI22_X1 U1155 ( .A1(n15023), .A2(n16017), .B1(n14699), .B2(n15021), .ZN(
        n1916) );
  OAI22_X1 U1156 ( .A1(n15022), .A2(n16016), .B1(n14702), .B2(n15020), .ZN(
        n1917) );
  OAI22_X1 U1157 ( .A1(n15131), .A2(n16015), .B1(n14669), .B2(n15127), .ZN(
        n1682) );
  OAI22_X1 U1158 ( .A1(n15131), .A2(n16014), .B1(n14690), .B2(n15127), .ZN(
        n1689) );
  OAI22_X1 U1159 ( .A1(n15128), .A2(n15979), .B1(n14633), .B2(n15126), .ZN(
        n3438) );
  OAI22_X1 U1160 ( .A1(n15129), .A2(n15978), .B1(n14640), .B2(n15126), .ZN(
        n3436) );
  OAI22_X1 U1161 ( .A1(n15133), .A2(n15977), .B1(n14651), .B2(n15126), .ZN(
        n1676) );
  OAI22_X1 U1162 ( .A1(n15129), .A2(n15976), .B1(n14673), .B2(n15126), .ZN(
        n3435) );
  OAI22_X1 U1163 ( .A1(n15130), .A2(n15974), .B1(n14702), .B2(n15127), .ZN(
        n1693) );
  OAI22_X1 U1164 ( .A1(n15131), .A2(n15961), .B1(n14681), .B2(n15127), .ZN(
        n1686) );
  OAI22_X1 U1165 ( .A1(n15027), .A2(n15947), .B1(n14633), .B2(n15020), .ZN(
        n1894) );
  OAI22_X1 U1166 ( .A1(n15027), .A2(n15945), .B1(n14639), .B2(n15020), .ZN(
        n1896) );
  OAI22_X1 U1167 ( .A1(n15026), .A2(n15944), .B1(n14648), .B2(n15020), .ZN(
        n1899) );
  OAI22_X1 U1168 ( .A1(n15026), .A2(n15926), .B1(n14642), .B2(n15020), .ZN(
        n1897) );
  OAI22_X1 U1169 ( .A1(n15045), .A2(n15918), .B1(n14669), .B2(n15040), .ZN(
        n2034) );
  OAI22_X1 U1170 ( .A1(n15043), .A2(n15917), .B1(n14690), .B2(n1110), .ZN(
        n2041) );
  OAI22_X1 U1171 ( .A1(n15048), .A2(n15912), .B1(n14625), .B2(n1110), .ZN(
        n2019) );
  OAI22_X1 U1172 ( .A1(n15168), .A2(n15886), .B1(n14704), .B2(n1087), .ZN(
        n1246) );
  OAI22_X1 U1173 ( .A1(n15228), .A2(n15865), .B1(n1082), .B2(n14659), .ZN(
        n1743) );
  OAI22_X1 U1174 ( .A1(n15197), .A2(n15864), .B1(n15204), .B2(n14707), .ZN(
        n1215) );
  OAI22_X1 U1175 ( .A1(n15160), .A2(n15806), .B1(n14647), .B2(n15153), .ZN(
        n1451) );
  OAI22_X1 U1176 ( .A1(n15159), .A2(n15798), .B1(n14662), .B2(n15153), .ZN(
        n1456) );
  OAI22_X1 U1177 ( .A1(n15166), .A2(n15910), .B1(n14668), .B2(n1087), .ZN(
        n3740) );
  OAI22_X1 U1178 ( .A1(n15167), .A2(n15908), .B1(n14689), .B2(n1087), .ZN(
        n3738) );
  OAI22_X1 U1179 ( .A1(n15172), .A2(n15891), .B1(n14620), .B2(n1087), .ZN(
        n1218) );
  OAI22_X1 U1180 ( .A1(n15171), .A2(n15890), .B1(n14635), .B2(n1087), .ZN(
        n1223) );
  OAI22_X1 U1181 ( .A1(n15170), .A2(n15889), .B1(n14674), .B2(n1087), .ZN(
        n1236) );
  OAI22_X1 U1182 ( .A1(n15169), .A2(n15887), .B1(n14692), .B2(n1087), .ZN(
        n1242) );
  OAI22_X1 U1183 ( .A1(n15096), .A2(n15854), .B1(n14664), .B2(n15088), .ZN(
        n3589) );
  OAI22_X1 U1184 ( .A1(n15227), .A2(n15842), .B1(n1082), .B2(n14671), .ZN(
        n1747) );
  OAI22_X1 U1185 ( .A1(n15077), .A2(n15841), .B1(n1097), .B2(n14623), .ZN(
        n1827) );
  OAI22_X1 U1186 ( .A1(n15077), .A2(n15840), .B1(n14630), .B2(n1097), .ZN(
        n1829) );
  OAI22_X1 U1187 ( .A1(n14984), .A2(n15582), .B1(n14662), .B2(n1123), .ZN(
        n1552) );
  OAI22_X1 U1188 ( .A1(n14963), .A2(n15504), .B1(n14662), .B2(n1125), .ZN(
        n1488) );
  OAI22_X1 U1189 ( .A1(n14959), .A2(n15498), .B1(n14712), .B2(n1125), .ZN(
        n1504) );
  OAI22_X1 U1190 ( .A1(n14963), .A2(n15432), .B1(n14660), .B2(n1125), .ZN(
        n1487) );
  OAI22_X1 U1191 ( .A1(n15048), .A2(n15789), .B1(n14630), .B2(n1110), .ZN(
        n2021) );
  OAI22_X1 U1192 ( .A1(n14995), .A2(n15749), .B1(n14669), .B2(n14990), .ZN(
        n1586) );
  OAI22_X1 U1193 ( .A1(n14993), .A2(n15748), .B1(n14690), .B2(n1122), .ZN(
        n1593) );
  OAI22_X1 U1194 ( .A1(n15230), .A2(n15723), .B1(n15222), .B2(n14632), .ZN(
        n1734) );
  OAI22_X1 U1195 ( .A1(n15229), .A2(n15722), .B1(n1082), .B2(n14638), .ZN(
        n1736) );
  OAI22_X1 U1196 ( .A1(n15110), .A2(n16205), .B1(n14621), .B2(n15108), .ZN(
        n3430) );
  OAI22_X1 U1197 ( .A1(n15110), .A2(n16204), .B1(n14636), .B2(n15108), .ZN(
        n3427) );
  OAI22_X1 U1198 ( .A1(n15111), .A2(n16203), .B1(n14675), .B2(n15108), .ZN(
        n3423) );
  OAI22_X1 U1199 ( .A1(n15111), .A2(n16202), .B1(n14687), .B2(n15108), .ZN(
        n3422) );
  OAI22_X1 U1200 ( .A1(n14961), .A2(n15680), .B1(n14686), .B2(n14958), .ZN(
        n1496) );
  OAI22_X1 U1201 ( .A1(n15160), .A2(n15701), .B1(n14646), .B2(n1088), .ZN(
        n1450) );
  OAI22_X1 U1202 ( .A1(n14965), .A2(n15580), .B1(n14643), .B2(n1125), .ZN(
        n1481) );
  OAI22_X1 U1203 ( .A1(n14987), .A2(n15530), .B1(n14621), .B2(n1123), .ZN(
        n1538) );
  OAI22_X1 U1204 ( .A1(n14986), .A2(n15529), .B1(n14636), .B2(n1123), .ZN(
        n1543) );
  OAI22_X1 U1205 ( .A1(n14982), .A2(n15525), .B1(n14687), .B2(n1123), .ZN(
        n1560) );
  OAI22_X1 U1206 ( .A1(n15112), .A2(n16292), .B1(n14711), .B2(n15109), .ZN(
        n1728) );
  OAI22_X1 U1207 ( .A1(n15112), .A2(n16291), .B1(n14714), .B2(n15109), .ZN(
        n1729) );
  OAI22_X1 U1208 ( .A1(n15025), .A2(n16163), .B1(n14660), .B2(n15021), .ZN(
        n1903) );
  OAI22_X1 U1209 ( .A1(n15169), .A2(n15888), .B1(n14686), .B2(n1087), .ZN(
        n1240) );
  OAI22_X1 U1210 ( .A1(n15114), .A2(n16265), .B1(n14669), .B2(n15109), .ZN(
        n1714) );
  OAI22_X1 U1211 ( .A1(n15140), .A2(n16256), .B1(n14669), .B2(n15136), .ZN(
        n3448) );
  OAI22_X1 U1212 ( .A1(n15141), .A2(n16255), .B1(n14690), .B2(n15136), .ZN(
        n3444) );
  OAI22_X1 U1213 ( .A1(n15238), .A2(n16239), .B1(n1081), .B2(n14665), .ZN(
        n3477) );
  OAI22_X1 U1214 ( .A1(n15238), .A2(n16238), .B1(n1081), .B2(n14677), .ZN(
        n3476) );
  OAI22_X1 U1215 ( .A1(n15239), .A2(n16237), .B1(n15233), .B2(n14695), .ZN(
        n3473) );
  OAI22_X1 U1216 ( .A1(n15124), .A2(n16218), .B1(n14653), .B2(n15117), .ZN(
        n1325) );
  OAI22_X1 U1217 ( .A1(n15124), .A2(n16217), .B1(n14656), .B2(n15118), .ZN(
        n1326) );
  OAI22_X1 U1218 ( .A1(n15119), .A2(n16216), .B1(n14680), .B2(n15117), .ZN(
        n3607) );
  OAI22_X1 U1219 ( .A1(n15123), .A2(n16215), .B1(n14683), .B2(n15118), .ZN(
        n1335) );
  OAI22_X1 U1220 ( .A1(n15115), .A2(n16194), .B1(n14654), .B2(n15108), .ZN(
        n1709) );
  OAI22_X1 U1221 ( .A1(n15114), .A2(n16193), .B1(n14657), .B2(n15109), .ZN(
        n1710) );
  OAI22_X1 U1222 ( .A1(n15247), .A2(n16150), .B1(n15254), .B2(n14641), .ZN(
        n2057) );
  OAI22_X1 U1223 ( .A1(n15130), .A2(n15975), .B1(n14699), .B2(n15127), .ZN(
        n1692) );
  OAI22_X1 U1224 ( .A1(n15058), .A2(n16128), .B1(n14649), .B2(n15051), .ZN(
        n3390) );
  OAI22_X1 U1225 ( .A1(n15059), .A2(n15990), .B1(n14685), .B2(n15051), .ZN(
        n2103) );
  OAI22_X1 U1226 ( .A1(n15134), .A2(n15980), .B1(n14627), .B2(n15127), .ZN(
        n1668) );
  OAI22_X1 U1227 ( .A1(n15170), .A2(n15909), .B1(n14671), .B2(n15164), .ZN(
        n1235) );
  OAI22_X1 U1228 ( .A1(n15048), .A2(n15903), .B1(n14633), .B2(n1110), .ZN(
        n2022) );
  OAI22_X1 U1229 ( .A1(n15047), .A2(n15901), .B1(n14639), .B2(n1110), .ZN(
        n2024) );
  OAI22_X1 U1230 ( .A1(n15046), .A2(n15898), .B1(n14663), .B2(n1110), .ZN(
        n2032) );
  OAI22_X1 U1231 ( .A1(n15044), .A2(n15896), .B1(n14675), .B2(n1110), .ZN(
        n2036) );
  OAI22_X1 U1232 ( .A1(n15045), .A2(n15895), .B1(n14687), .B2(n1110), .ZN(
        n2040) );
  OAI22_X1 U1233 ( .A1(n15043), .A2(n15894), .B1(n14693), .B2(n1110), .ZN(
        n2042) );
  OAI22_X1 U1234 ( .A1(n15044), .A2(n15893), .B1(n14705), .B2(n1110), .ZN(
        n2046) );
  OAI22_X1 U1235 ( .A1(n15167), .A2(n15850), .B1(n1087), .B2(n14707), .ZN(
        n1247) );
  OAI22_X1 U1236 ( .A1(n15167), .A2(n15818), .B1(n1087), .B2(n14710), .ZN(
        n1248) );
  OAI22_X1 U1237 ( .A1(n15167), .A2(n15817), .B1(n1087), .B2(n14713), .ZN(
        n1249) );
  OAI22_X1 U1238 ( .A1(n15166), .A2(n15768), .B1(n14664), .B2(n1087), .ZN(
        n3741) );
  OAI22_X1 U1239 ( .A1(n15096), .A2(n15714), .B1(n1095), .B2(n14624), .ZN(
        n1155) );
  OAI22_X1 U1240 ( .A1(n15158), .A2(n15700), .B1(n14671), .B2(n15153), .ZN(
        n1459) );
  OAI22_X1 U1241 ( .A1(n15156), .A2(n15699), .B1(n1088), .B2(n14707), .ZN(
        n3730) );
  OAI22_X1 U1242 ( .A1(n15161), .A2(n15696), .B1(n14632), .B2(n1088), .ZN(
        n1446) );
  OAI22_X1 U1243 ( .A1(n15160), .A2(n15695), .B1(n14638), .B2(n1088), .ZN(
        n1448) );
  OAI22_X1 U1244 ( .A1(n15159), .A2(n15694), .B1(n14661), .B2(n1088), .ZN(
        n1455) );
  OAI22_X1 U1245 ( .A1(n14984), .A2(n15528), .B1(n14666), .B2(n1123), .ZN(
        n1553) );
  OAI22_X1 U1246 ( .A1(n14983), .A2(n15527), .B1(n14675), .B2(n14979), .ZN(
        n1556) );
  OAI22_X1 U1247 ( .A1(n14983), .A2(n15526), .B1(n14678), .B2(n1123), .ZN(
        n1557) );
  OAI22_X1 U1248 ( .A1(n14982), .A2(n15524), .B1(n14693), .B2(n1123), .ZN(
        n1562) );
  OAI22_X1 U1249 ( .A1(n14982), .A2(n15523), .B1(n14696), .B2(n1123), .ZN(
        n1563) );
  OAI22_X1 U1250 ( .A1(n14981), .A2(n15522), .B1(n14705), .B2(n1123), .ZN(
        n1566) );
  OAI22_X1 U1251 ( .A1(n14981), .A2(n15510), .B1(n14709), .B2(n14979), .ZN(
        n1567) );
  OAI22_X1 U1252 ( .A1(n14962), .A2(n15509), .B1(n14671), .B2(n14958), .ZN(
        n1491) );
  OAI22_X1 U1253 ( .A1(n14987), .A2(n15503), .B1(n14627), .B2(n14979), .ZN(
        n1540) );
  OAI22_X1 U1254 ( .A1(n14985), .A2(n15502), .B1(n14651), .B2(n14979), .ZN(
        n1548) );
  OAI22_X1 U1255 ( .A1(n14981), .A2(n15500), .B1(n14702), .B2(n1123), .ZN(
        n1565) );
  OAI22_X1 U1256 ( .A1(n15138), .A2(n16303), .B1(n14707), .B2(n15135), .ZN(
        n3614) );
  OAI22_X1 U1257 ( .A1(n15113), .A2(n16264), .B1(n14690), .B2(n15109), .ZN(
        n1721) );
  OAI22_X1 U1258 ( .A1(n15110), .A2(n16192), .B1(n14680), .B2(n15109), .ZN(
        n3606) );
  OAI22_X1 U1259 ( .A1(n15113), .A2(n16191), .B1(n14684), .B2(n15109), .ZN(
        n1719) );
  OAI22_X1 U1260 ( .A1(n15114), .A2(n16184), .B1(n14660), .B2(n15109), .ZN(
        n1711) );
  OAI22_X1 U1261 ( .A1(n15055), .A2(n16170), .B1(n14629), .B2(n15050), .ZN(
        n3509) );
  OAI22_X1 U1262 ( .A1(n15129), .A2(n16093), .B1(n14675), .B2(n15126), .ZN(
        n3434) );
  OAI22_X1 U1263 ( .A1(n15129), .A2(n16092), .B1(n14687), .B2(n15126), .ZN(
        n3433) );
  OAI22_X1 U1264 ( .A1(n15054), .A2(n16052), .B1(n14644), .B2(n15050), .ZN(
        n3506) );
  OAI22_X1 U1265 ( .A1(n15027), .A2(n16022), .B1(n14630), .B2(n15020), .ZN(
        n1893) );
  OAI22_X1 U1266 ( .A1(n15025), .A2(n16020), .B1(n14666), .B2(n15021), .ZN(
        n1905) );
  OAI22_X1 U1267 ( .A1(n15024), .A2(n16019), .B1(n14678), .B2(n15021), .ZN(
        n1909) );
  OAI22_X1 U1268 ( .A1(n15053), .A2(n16007), .B1(n14626), .B2(n15050), .ZN(
        n3510) );
  OAI22_X1 U1269 ( .A1(n15054), .A2(n16006), .B1(n14650), .B2(n15050), .ZN(
        n3505) );
  OAI22_X1 U1270 ( .A1(n15055), .A2(n16004), .B1(n14666), .B2(n15050), .ZN(
        n3503) );
  OAI22_X1 U1271 ( .A1(n15056), .A2(n16003), .B1(n14677), .B2(n15050), .ZN(
        n3500) );
  OAI22_X1 U1272 ( .A1(n15056), .A2(n16002), .B1(n14696), .B2(n15051), .ZN(
        n3498) );
  OAI22_X1 U1273 ( .A1(n15056), .A2(n16001), .B1(n14698), .B2(n15051), .ZN(
        n3497) );
  OAI22_X1 U1274 ( .A1(n15057), .A2(n16000), .B1(n14702), .B2(n15051), .ZN(
        n3496) );
  OAI22_X1 U1275 ( .A1(n15059), .A2(n15993), .B1(n14655), .B2(n15051), .ZN(
        n2093) );
  OAI22_X1 U1276 ( .A1(n15059), .A2(n15992), .B1(n14658), .B2(n15051), .ZN(
        n2094) );
  OAI22_X1 U1277 ( .A1(n15059), .A2(n15991), .B1(n14680), .B2(n15051), .ZN(
        n2102) );
  OAI22_X1 U1278 ( .A1(n15133), .A2(n15954), .B1(n14642), .B2(n15126), .ZN(
        n1673) );
  OAI22_X1 U1279 ( .A1(n15133), .A2(n15953), .B1(n14645), .B2(n15127), .ZN(
        n1674) );
  OAI22_X1 U1280 ( .A1(n15026), .A2(n15925), .B1(n14645), .B2(n15020), .ZN(
        n1898) );
  OAI22_X1 U1281 ( .A1(n15067), .A2(n15958), .B1(n14657), .B2(n15060), .ZN(
        n1870) );
  OAI22_X1 U1282 ( .A1(n15048), .A2(n15904), .B1(n14621), .B2(n1110), .ZN(
        n2018) );
  OAI22_X1 U1283 ( .A1(n15045), .A2(n15902), .B1(n14636), .B2(n15040), .ZN(
        n2023) );
  OAI22_X1 U1284 ( .A1(n15158), .A2(n15863), .B1(n14641), .B2(n1088), .ZN(
        n3734) );
  OAI22_X1 U1285 ( .A1(n15166), .A2(n15851), .B1(n14659), .B2(n1087), .ZN(
        n3742) );
  OAI22_X1 U1286 ( .A1(n15198), .A2(n15816), .B1(n15205), .B2(n14680), .ZN(
        n1206) );
  OAI22_X1 U1287 ( .A1(n14986), .A2(n15670), .B1(n14642), .B2(n1123), .ZN(
        n1545) );
  OAI22_X1 U1288 ( .A1(n14986), .A2(n15669), .B1(n14645), .B2(n1123), .ZN(
        n1546) );
  OAI22_X1 U1289 ( .A1(n14996), .A2(n15645), .B1(n14661), .B2(n1122), .ZN(
        n1583) );
  OAI22_X1 U1290 ( .A1(n15004), .A2(n15780), .B1(n14681), .B2(n15001), .ZN(
        n1622) );
  OAI22_X1 U1291 ( .A1(n14997), .A2(n15731), .B1(n14642), .B2(n1122), .ZN(
        n1577) );
  OAI22_X1 U1292 ( .A1(n14985), .A2(n15513), .B1(n14653), .B2(n14979), .ZN(
        n1549) );
  OAI22_X1 U1293 ( .A1(n14985), .A2(n15512), .B1(n14656), .B2(n1123), .ZN(
        n1550) );
  OAI22_X1 U1294 ( .A1(n14981), .A2(n15501), .B1(n14699), .B2(n1123), .ZN(
        n1564) );
  OAI22_X1 U1295 ( .A1(n15132), .A2(n16127), .B1(n14654), .B2(n15126), .ZN(
        n1677) );
  OAI22_X1 U1296 ( .A1(n15132), .A2(n16126), .B1(n14657), .B2(n15127), .ZN(
        n1678) );
  OAI22_X1 U1297 ( .A1(n15131), .A2(n16125), .B1(n14684), .B2(n15127), .ZN(
        n1687) );
  OAI22_X1 U1298 ( .A1(n15130), .A2(n16124), .B1(n14708), .B2(n15126), .ZN(
        n1695) );
  OAI22_X1 U1299 ( .A1(n15128), .A2(n16096), .B1(n14621), .B2(n15126), .ZN(
        n3439) );
  OAI22_X1 U1300 ( .A1(n15128), .A2(n16094), .B1(n14636), .B2(n15126), .ZN(
        n3437) );
  OAI22_X1 U1301 ( .A1(n15129), .A2(n16091), .B1(n14693), .B2(n15126), .ZN(
        n3432) );
  OAI22_X1 U1302 ( .A1(n15130), .A2(n16090), .B1(n14705), .B2(n15126), .ZN(
        n3431) );
  OAI22_X1 U1303 ( .A1(n15125), .A2(n16086), .B1(n14632), .B2(n15117), .ZN(
        n1318) );
  OAI22_X1 U1304 ( .A1(n15124), .A2(n16085), .B1(n14638), .B2(n15118), .ZN(
        n1320) );
  OAI22_X1 U1305 ( .A1(n15081), .A2(n16121), .B1(n14677), .B2(n15080), .ZN(
        n3581) );
  OAI22_X1 U1306 ( .A1(n15083), .A2(n16075), .B1(n14655), .B2(n15079), .ZN(
        n3407) );
  OAI22_X1 U1307 ( .A1(n15083), .A2(n16074), .B1(n14658), .B2(n15080), .ZN(
        n3406) );
  OAI22_X1 U1308 ( .A1(n15084), .A2(n16073), .B1(n14685), .B2(n15080), .ZN(
        n3400) );
  OAI22_X1 U1309 ( .A1(n15086), .A2(n16072), .B1(n14708), .B2(n15080), .ZN(
        n1791) );
  OAI22_X1 U1310 ( .A1(n15066), .A2(n16039), .B1(n14708), .B2(n15061), .ZN(
        n1887) );
  OAI22_X1 U1311 ( .A1(n15105), .A2(n16032), .B1(n14670), .B2(n15100), .ZN(
        n1266) );
  OAI22_X1 U1312 ( .A1(n15104), .A2(n16031), .B1(n14691), .B2(n15100), .ZN(
        n1273) );
  OAI22_X1 U1313 ( .A1(n15084), .A2(n16025), .B1(n14681), .B2(n15080), .ZN(
        n3401) );
  OAI22_X1 U1314 ( .A1(n15023), .A2(n16018), .B1(n14696), .B2(n15021), .ZN(
        n1915) );
  OAI22_X1 U1315 ( .A1(n15067), .A2(n15959), .B1(n14654), .B2(n15061), .ZN(
        n1869) );
  OAI22_X1 U1316 ( .A1(n15067), .A2(n15957), .B1(n14681), .B2(n15060), .ZN(
        n1878) );
  OAI22_X1 U1317 ( .A1(n15066), .A2(n15956), .B1(n14684), .B2(n15061), .ZN(
        n1879) );
  OAI22_X1 U1318 ( .A1(n15132), .A2(n15931), .B1(n14663), .B2(n15127), .ZN(
        n1680) );
  OAI22_X1 U1319 ( .A1(n15022), .A2(n15924), .B1(n14711), .B2(n15020), .ZN(
        n1920) );
  OAI22_X1 U1320 ( .A1(n15022), .A2(n15923), .B1(n14714), .B2(n15021), .ZN(
        n1921) );
  OAI22_X1 U1321 ( .A1(n15047), .A2(n15900), .B1(n14648), .B2(n15040), .ZN(
        n2027) );
  OAI22_X1 U1322 ( .A1(n15045), .A2(n15897), .B1(n14672), .B2(n1110), .ZN(
        n2035) );
  OAI22_X1 U1323 ( .A1(n15081), .A2(n15930), .B1(n14627), .B2(n15079), .ZN(
        n3416) );
  OAI22_X1 U1324 ( .A1(n15085), .A2(n15928), .B1(n14699), .B2(n15080), .ZN(
        n3396) );
  OAI22_X1 U1325 ( .A1(n15172), .A2(n15852), .B1(n1087), .B2(n14624), .ZN(
        n1219) );
  OAI22_X1 U1326 ( .A1(n15156), .A2(n15844), .B1(n1088), .B2(n14710), .ZN(
        n1472) );
  OAI22_X1 U1327 ( .A1(n15157), .A2(n15843), .B1(n1088), .B2(n14713), .ZN(
        n1473) );
  OAI22_X1 U1328 ( .A1(n15172), .A2(n15832), .B1(n14628), .B2(n1087), .ZN(
        n1220) );
  OAI22_X1 U1329 ( .A1(n15172), .A2(n15831), .B1(n14631), .B2(n15164), .ZN(
        n1221) );
  OAI22_X1 U1330 ( .A1(n15171), .A2(n15829), .B1(n14646), .B2(n15164), .ZN(
        n1226) );
  OAI22_X1 U1331 ( .A1(n15171), .A2(n15828), .B1(n14652), .B2(n1087), .ZN(
        n1228) );
  OAI22_X1 U1332 ( .A1(n15170), .A2(n15827), .B1(n14667), .B2(n1087), .ZN(
        n1233) );
  OAI22_X1 U1333 ( .A1(n15170), .A2(n15826), .B1(n14679), .B2(n1087), .ZN(
        n1237) );
  OAI22_X1 U1334 ( .A1(n15168), .A2(n15825), .B1(n14697), .B2(n1087), .ZN(
        n1243) );
  OAI22_X1 U1335 ( .A1(n15168), .A2(n15824), .B1(n14700), .B2(n15164), .ZN(
        n1244) );
  OAI22_X1 U1336 ( .A1(n15168), .A2(n15823), .B1(n14703), .B2(n1087), .ZN(
        n1245) );
  OAI22_X1 U1337 ( .A1(n15047), .A2(n15788), .B1(n14641), .B2(n15040), .ZN(
        n2025) );
  OAI22_X1 U1338 ( .A1(n15047), .A2(n15787), .B1(n14644), .B2(n15040), .ZN(
        n2026) );
  OAI22_X1 U1339 ( .A1(n14976), .A2(n15775), .B1(n14624), .B2(n1124), .ZN(
        n1507) );
  OAI22_X1 U1340 ( .A1(n14974), .A2(n15774), .B1(n14661), .B2(n1124), .ZN(
        n1519) );
  OAI22_X1 U1341 ( .A1(n15171), .A2(n15771), .B1(n14632), .B2(n15164), .ZN(
        n3747) );
  OAI22_X1 U1342 ( .A1(n15165), .A2(n15770), .B1(n14638), .B2(n1087), .ZN(
        n3746) );
  OAI22_X1 U1343 ( .A1(n15166), .A2(n15769), .B1(n14647), .B2(n1087), .ZN(
        n3745) );
  OAI22_X1 U1344 ( .A1(n14975), .A2(n15766), .B1(n14642), .B2(n1124), .ZN(
        n1513) );
  OAI22_X1 U1345 ( .A1(n14974), .A2(n15765), .B1(n14645), .B2(n1124), .ZN(
        n1514) );
  OAI22_X1 U1346 ( .A1(n15159), .A2(n15725), .B1(n14670), .B2(n15153), .ZN(
        n1458) );
  OAI22_X1 U1347 ( .A1(n15157), .A2(n15724), .B1(n14691), .B2(n1088), .ZN(
        n1465) );
  OAI22_X1 U1348 ( .A1(n15180), .A2(n15715), .B1(n14663), .B2(n1086), .ZN(
        n1968) );
  OAI22_X1 U1349 ( .A1(n14983), .A2(n15585), .B1(n14681), .B2(n1123), .ZN(
        n1558) );
  OAI22_X1 U1350 ( .A1(n14987), .A2(n15579), .B1(n14624), .B2(n14979), .ZN(
        n1539) );
  OAI22_X1 U1351 ( .A1(n14983), .A2(n15511), .B1(n14683), .B2(n1123), .ZN(
        n1559) );
  OAI22_X1 U1352 ( .A1(n15161), .A2(n15666), .B1(n14628), .B2(n15153), .ZN(
        n1444) );
  OAI22_X1 U1353 ( .A1(n15157), .A2(n15659), .B1(n14703), .B2(n1088), .ZN(
        n1469) );
  OAI22_X1 U1354 ( .A1(n14985), .A2(n15581), .B1(n14661), .B2(n1123), .ZN(
        n1551) );
  OAI22_X1 U1355 ( .A1(n15005), .A2(n15540), .B1(n14669), .B2(n15001), .ZN(
        n1618) );
  OAI22_X1 U1356 ( .A1(n15003), .A2(n15539), .B1(n14690), .B2(n15001), .ZN(
        n1625) );
  OAI22_X1 U1357 ( .A1(n14980), .A2(n15521), .B1(n14712), .B2(n1123), .ZN(
        n1568) );
  OAI22_X1 U1358 ( .A1(n14984), .A2(n15520), .B1(n14715), .B2(n1123), .ZN(
        n1569) );
  OAI22_X1 U1359 ( .A1(n15006), .A2(n15437), .B1(n14654), .B2(n15000), .ZN(
        n1613) );
  OAI22_X1 U1360 ( .A1(n15005), .A2(n15436), .B1(n14657), .B2(n15001), .ZN(
        n1614) );
  OAI22_X1 U1361 ( .A1(n15004), .A2(n15435), .B1(n14684), .B2(n15001), .ZN(
        n1623) );
  OAI22_X1 U1362 ( .A1(n15106), .A2(n16166), .B1(n14653), .B2(n15100), .ZN(
        n1261) );
  OAI22_X1 U1363 ( .A1(n15106), .A2(n16165), .B1(n14656), .B2(n15099), .ZN(
        n1262) );
  OAI22_X1 U1364 ( .A1(n15104), .A2(n16164), .B1(n14683), .B2(n15100), .ZN(
        n1271) );
  OAI22_X1 U1365 ( .A1(n15104), .A2(n16139), .B1(n14708), .B2(n15100), .ZN(
        n3565) );
  OAI22_X1 U1366 ( .A1(n15081), .A2(n16123), .B1(n14630), .B2(n15079), .ZN(
        n3415) );
  OAI22_X1 U1367 ( .A1(n15084), .A2(n16122), .B1(n14665), .B2(n15080), .ZN(
        n3404) );
  OAI22_X1 U1368 ( .A1(n15085), .A2(n16120), .B1(n14695), .B2(n15080), .ZN(
        n3397) );
  OAI22_X1 U1369 ( .A1(n15063), .A2(n16088), .B1(n14644), .B2(n15060), .ZN(
        n3526) );
  OAI22_X1 U1370 ( .A1(n15161), .A2(n15667), .B1(n1088), .B2(n14624), .ZN(
        n1443) );
  OAI22_X1 U1371 ( .A1(n15105), .A2(n16067), .B1(n14682), .B2(n15100), .ZN(
        n1270) );
  OAI22_X1 U1372 ( .A1(n15025), .A2(n16064), .B1(n14669), .B2(n15021), .ZN(
        n1906) );
  OAI22_X1 U1373 ( .A1(n15087), .A2(n16026), .B1(n14669), .B2(n15079), .ZN(
        n1778) );
  OAI22_X1 U1374 ( .A1(n15086), .A2(n16024), .B1(n14690), .B2(n15080), .ZN(
        n1785) );
  OAI22_X1 U1375 ( .A1(n15081), .A2(n15955), .B1(n15080), .B2(n14623), .ZN(
        n3417) );
  OAI22_X1 U1376 ( .A1(n15065), .A2(n16013), .B1(n14711), .B2(n15061), .ZN(
        n3513) );
  OAI22_X1 U1377 ( .A1(n15065), .A2(n16012), .B1(n14714), .B2(n15061), .ZN(
        n3512) );
  OAI22_X1 U1378 ( .A1(n15083), .A2(n15929), .B1(n14651), .B2(n15079), .ZN(
        n3408) );
  OAI22_X1 U1379 ( .A1(n15085), .A2(n15927), .B1(n14702), .B2(n15079), .ZN(
        n3395) );
  OAI22_X1 U1380 ( .A1(n15169), .A2(n15905), .B1(n14682), .B2(n15164), .ZN(
        n1238) );
  OAI22_X1 U1381 ( .A1(n14976), .A2(n15713), .B1(n14621), .B2(n14968), .ZN(
        n1506) );
  OAI22_X1 U1382 ( .A1(n14975), .A2(n15711), .B1(n14636), .B2(n14968), .ZN(
        n1511) );
  OAI22_X1 U1383 ( .A1(n14972), .A2(n15707), .B1(n14671), .B2(n1124), .ZN(
        n1523) );
  OAI22_X1 U1384 ( .A1(n14972), .A2(n15706), .B1(n14675), .B2(n1124), .ZN(
        n1524) );
  OAI22_X1 U1385 ( .A1(n14971), .A2(n15704), .B1(n14693), .B2(n1124), .ZN(
        n1530) );
  OAI22_X1 U1386 ( .A1(n15161), .A2(n15665), .B1(n14631), .B2(n1088), .ZN(
        n1445) );
  OAI22_X1 U1387 ( .A1(n15158), .A2(n15662), .B1(n14679), .B2(n1088), .ZN(
        n1461) );
  OAI22_X1 U1388 ( .A1(n15157), .A2(n15661), .B1(n14697), .B2(n1088), .ZN(
        n1467) );
  OAI22_X1 U1389 ( .A1(n15158), .A2(n15660), .B1(n14700), .B2(n1088), .ZN(
        n1468) );
  OAI22_X1 U1390 ( .A1(n15004), .A2(n15628), .B1(n14672), .B2(n15001), .ZN(
        n1619) );
  OAI22_X1 U1391 ( .A1(n15023), .A2(n16061), .B1(n14690), .B2(n15021), .ZN(
        n1913) );
  OAI22_X1 U1392 ( .A1(n15028), .A2(n15921), .B1(n14625), .B2(n15020), .ZN(
        n1891) );
  OAI22_X1 U1393 ( .A1(n14976), .A2(n15779), .B1(n14628), .B2(n1124), .ZN(
        n1508) );
  OAI22_X1 U1394 ( .A1(n14970), .A2(n15777), .B1(n14700), .B2(n14968), .ZN(
        n1532) );
  OAI22_X1 U1395 ( .A1(n14972), .A2(n15705), .B1(n14687), .B2(n1124), .ZN(
        n1528) );
  OAI22_X1 U1396 ( .A1(n14970), .A2(n15703), .B1(n14705), .B2(n1124), .ZN(
        n1534) );
  OAI22_X1 U1397 ( .A1(n14970), .A2(n15702), .B1(n14709), .B2(n1124), .ZN(
        n1535) );
  OAI22_X1 U1398 ( .A1(n15160), .A2(n15664), .B1(n14652), .B2(n1088), .ZN(
        n1452) );
  OAI22_X1 U1399 ( .A1(n15159), .A2(n15663), .B1(n14667), .B2(n15153), .ZN(
        n1457) );
  OAI22_X1 U1400 ( .A1(n15007), .A2(n15741), .B1(n14633), .B2(n15000), .ZN(
        n1606) );
  OAI22_X1 U1401 ( .A1(n15007), .A2(n15740), .B1(n14639), .B2(n15000), .ZN(
        n1608) );
  OAI22_X1 U1402 ( .A1(n15014), .A2(n15560), .B1(n14663), .B2(n1119), .ZN(
        n1808) );
  OAI22_X1 U1403 ( .A1(n15212), .A2(n15495), .B1(n15218), .B2(n14689), .ZN(
        n1401) );
  OAI22_X1 U1404 ( .A1(n15101), .A2(n16147), .B1(n14620), .B2(n15099), .ZN(
        n3605) );
  OAI22_X1 U1405 ( .A1(n15101), .A2(n16146), .B1(n14635), .B2(n15099), .ZN(
        n3604) );
  OAI22_X1 U1406 ( .A1(n15105), .A2(n16145), .B1(n14671), .B2(n15100), .ZN(
        n1267) );
  OAI22_X1 U1407 ( .A1(n15101), .A2(n16144), .B1(n14674), .B2(n15099), .ZN(
        n3603) );
  OAI22_X1 U1408 ( .A1(n15101), .A2(n16143), .B1(n14686), .B2(n15099), .ZN(
        n3602) );
  OAI22_X1 U1409 ( .A1(n15101), .A2(n16142), .B1(n14692), .B2(n15099), .ZN(
        n3601) );
  OAI22_X1 U1410 ( .A1(n15102), .A2(n16141), .B1(n14704), .B2(n15099), .ZN(
        n3600) );
  OAI22_X1 U1411 ( .A1(n15081), .A2(n16138), .B1(n14621), .B2(n15079), .ZN(
        n3418) );
  OAI22_X1 U1412 ( .A1(n15084), .A2(n16136), .B1(n14672), .B2(n15080), .ZN(
        n3403) );
  OAI22_X1 U1413 ( .A1(n15084), .A2(n16135), .B1(n14675), .B2(n15080), .ZN(
        n3402) );
  OAI22_X1 U1414 ( .A1(n15085), .A2(n16134), .B1(n14687), .B2(n15080), .ZN(
        n3399) );
  OAI22_X1 U1415 ( .A1(n15085), .A2(n16133), .B1(n14693), .B2(n15080), .ZN(
        n3398) );
  OAI22_X1 U1416 ( .A1(n15086), .A2(n16132), .B1(n14705), .B2(n15079), .ZN(
        n3394) );
  OAI22_X1 U1417 ( .A1(n15015), .A2(n15729), .B1(n14660), .B2(n15009), .ZN(
        n1807) );
  OAI22_X1 U1418 ( .A1(n15062), .A2(n16117), .B1(n14629), .B2(n15060), .ZN(
        n3530) );
  OAI22_X1 U1419 ( .A1(n15063), .A2(n16115), .B1(n14651), .B2(n15060), .ZN(
        n3524) );
  OAI22_X1 U1420 ( .A1(n15064), .A2(n16113), .B1(n14673), .B2(n15061), .ZN(
        n3519) );
  OAI22_X1 U1421 ( .A1(n15064), .A2(n16111), .B1(n14677), .B2(n15061), .ZN(
        n3518) );
  OAI22_X1 U1422 ( .A1(n15102), .A2(n16083), .B1(n14626), .B2(n15099), .ZN(
        n3574) );
  OAI22_X1 U1423 ( .A1(n15103), .A2(n16077), .B1(n14698), .B2(n15100), .ZN(
        n3567) );
  OAI22_X1 U1424 ( .A1(n15103), .A2(n16076), .B1(n14701), .B2(n15100), .ZN(
        n3566) );
  OAI22_X1 U1425 ( .A1(n15106), .A2(n16069), .B1(n14647), .B2(n15099), .ZN(
        n1259) );
  OAI22_X1 U1426 ( .A1(n15068), .A2(n16045), .B1(n15061), .B2(n14623), .ZN(
        n1859) );
  OAI22_X1 U1427 ( .A1(n15063), .A2(n16042), .B1(n14649), .B2(n15060), .ZN(
        n3525) );
  OAI22_X1 U1428 ( .A1(n15082), .A2(n16029), .B1(n14639), .B2(n15079), .ZN(
        n3412) );
  OAI22_X1 U1429 ( .A1(n15102), .A2(n15936), .B1(n14641), .B2(n15099), .ZN(
        n3573) );
  OAI22_X1 U1430 ( .A1(n15102), .A2(n15935), .B1(n14644), .B2(n15099), .ZN(
        n3572) );
  OAI22_X1 U1431 ( .A1(n14971), .A2(n15919), .B1(n14691), .B2(n1124), .ZN(
        n1529) );
  OAI22_X1 U1432 ( .A1(n14971), .A2(n15833), .B1(n14681), .B2(n1124), .ZN(
        n1526) );
  OAI22_X1 U1433 ( .A1(n14974), .A2(n15778), .B1(n14652), .B2(n1124), .ZN(
        n1516) );
  OAI22_X1 U1434 ( .A1(n14970), .A2(n15776), .B1(n14703), .B2(n1124), .ZN(
        n1533) );
  OAI22_X1 U1435 ( .A1(n15212), .A2(n15496), .B1(n15219), .B2(n14668), .ZN(
        n1394) );
  OAI22_X1 U1436 ( .A1(n15008), .A2(n15747), .B1(n14625), .B2(n15000), .ZN(
        n1603) );
  OAI22_X1 U1437 ( .A1(n15005), .A2(n15746), .B1(n14660), .B2(n15001), .ZN(
        n1615) );
  OAI22_X1 U1438 ( .A1(n15189), .A2(n15744), .B1(n14657), .B2(n1085), .ZN(
        n1934) );
  OAI22_X1 U1439 ( .A1(n15188), .A2(n15743), .B1(n14684), .B2(n1085), .ZN(
        n1943) );
  OAI22_X1 U1440 ( .A1(n15186), .A2(n15742), .B1(n15184), .B2(n14707), .ZN(
        n1951) );
  OAI22_X1 U1441 ( .A1(n15006), .A2(n15739), .B1(n14648), .B2(n15000), .ZN(
        n1611) );
  OAI22_X1 U1442 ( .A1(n15005), .A2(n15738), .B1(n14662), .B2(n15001), .ZN(
        n1616) );
  OAI22_X1 U1443 ( .A1(n15211), .A2(n15734), .B1(n14653), .B2(n15214), .ZN(
        n1389) );
  OAI22_X1 U1444 ( .A1(n15212), .A2(n15733), .B1(n14656), .B2(n15213), .ZN(
        n1390) );
  OAI22_X1 U1445 ( .A1(n15212), .A2(n15732), .B1(n14683), .B2(n15214), .ZN(
        n1399) );
  OAI22_X1 U1446 ( .A1(n15017), .A2(n15730), .B1(n14625), .B2(n1119), .ZN(
        n1795) );
  OAI22_X1 U1447 ( .A1(n15014), .A2(n15728), .B1(n14666), .B2(n1119), .ZN(
        n1809) );
  OAI22_X1 U1448 ( .A1(n15013), .A2(n15727), .B1(n14678), .B2(n1119), .ZN(
        n1813) );
  OAI22_X1 U1449 ( .A1(n15012), .A2(n15726), .B1(n14696), .B2(n1119), .ZN(
        n1819) );
  OAI22_X1 U1450 ( .A1(n15064), .A2(n16114), .B1(n14665), .B2(n15060), .ZN(
        n3521) );
  OAI22_X1 U1451 ( .A1(n15086), .A2(n16034), .B1(n14711), .B2(n15080), .ZN(
        n3393) );
  OAI22_X1 U1452 ( .A1(n14975), .A2(n15712), .B1(n14632), .B2(n14968), .ZN(
        n1510) );
  OAI22_X1 U1453 ( .A1(n14975), .A2(n15710), .B1(n14638), .B2(n14968), .ZN(
        n1512) );
  OAI22_X1 U1454 ( .A1(n14974), .A2(n15709), .B1(n14647), .B2(n14968), .ZN(
        n1515) );
  OAI22_X1 U1455 ( .A1(n14973), .A2(n15708), .B1(n14662), .B2(n1124), .ZN(
        n1520) );
  OAI22_X1 U1456 ( .A1(n15006), .A2(n15644), .B1(n14651), .B2(n15000), .ZN(
        n1612) );
  OAI22_X1 U1457 ( .A1(n15005), .A2(n15643), .B1(n14666), .B2(n15001), .ZN(
        n1617) );
  OAI22_X1 U1458 ( .A1(n15004), .A2(n15642), .B1(n14678), .B2(n15001), .ZN(
        n1621) );
  OAI22_X1 U1459 ( .A1(n15003), .A2(n15641), .B1(n14696), .B2(n15000), .ZN(
        n1627) );
  OAI22_X1 U1460 ( .A1(n15003), .A2(n15640), .B1(n14699), .B2(n15001), .ZN(
        n1628) );
  OAI22_X1 U1461 ( .A1(n15002), .A2(n15639), .B1(n14702), .B2(n15000), .ZN(
        n1629) );
  OAI22_X1 U1462 ( .A1(n15002), .A2(n15561), .B1(n14714), .B2(n15001), .ZN(
        n1633) );
  OAI22_X1 U1463 ( .A1(n15185), .A2(n15555), .B1(n14668), .B2(n1085), .ZN(
        n3776) );
  OAI22_X1 U1464 ( .A1(n15107), .A2(n16140), .B1(n15100), .B2(n14624), .ZN(
        n1251) );
  OAI22_X1 U1465 ( .A1(n15082), .A2(n16137), .B1(n14636), .B2(n15079), .ZN(
        n3413) );
  OAI22_X1 U1466 ( .A1(n15062), .A2(n16118), .B1(n14627), .B2(n15061), .ZN(
        n3531) );
  OAI22_X1 U1467 ( .A1(n15066), .A2(n16110), .B1(n14687), .B2(n15060), .ZN(
        n1880) );
  OAI22_X1 U1468 ( .A1(n15066), .A2(n16109), .B1(n14693), .B2(n15061), .ZN(
        n1882) );
  OAI22_X1 U1469 ( .A1(n15065), .A2(n16108), .B1(n14695), .B2(n15061), .ZN(
        n3516) );
  OAI22_X1 U1470 ( .A1(n15065), .A2(n16107), .B1(n14699), .B2(n15061), .ZN(
        n3515) );
  OAI22_X1 U1471 ( .A1(n15065), .A2(n16106), .B1(n14701), .B2(n15061), .ZN(
        n3514) );
  OAI22_X1 U1472 ( .A1(n15066), .A2(n16105), .B1(n14705), .B2(n15061), .ZN(
        n1886) );
  OAI22_X1 U1473 ( .A1(n15106), .A2(n16071), .B1(n14632), .B2(n15100), .ZN(
        n1254) );
  OAI22_X1 U1474 ( .A1(n15106), .A2(n16070), .B1(n14638), .B2(n15099), .ZN(
        n1256) );
  OAI22_X1 U1475 ( .A1(n15105), .A2(n16068), .B1(n14662), .B2(n15100), .ZN(
        n1264) );
  OAI22_X1 U1476 ( .A1(n15083), .A2(n16028), .B1(n14649), .B2(n15079), .ZN(
        n3409) );
  OAI22_X1 U1477 ( .A1(n15083), .A2(n16027), .B1(n14663), .B2(n15080), .ZN(
        n3405) );
  OAI22_X1 U1478 ( .A1(n14973), .A2(n15920), .B1(n14670), .B2(n1124), .ZN(
        n1522) );
  OAI22_X1 U1479 ( .A1(n15212), .A2(n15611), .B1(n15218), .B2(n14674), .ZN(
        n1396) );
  OAI22_X1 U1480 ( .A1(n15002), .A2(n15562), .B1(n14711), .B2(n15000), .ZN(
        n1632) );
  OAI22_X1 U1481 ( .A1(n15007), .A2(n15558), .B1(n14627), .B2(n15000), .ZN(
        n1604) );
  OAI22_X1 U1482 ( .A1(n15067), .A2(n16112), .B1(n14675), .B2(n15061), .ZN(
        n1876) );
  OAI22_X1 U1483 ( .A1(n15062), .A2(n16089), .B1(n14641), .B2(n15060), .ZN(
        n3527) );
  OAI22_X1 U1484 ( .A1(n15102), .A2(n16081), .B1(n14650), .B2(n15099), .ZN(
        n3571) );
  OAI22_X1 U1485 ( .A1(n15103), .A2(n16080), .B1(n14665), .B2(n15099), .ZN(
        n3570) );
  OAI22_X1 U1486 ( .A1(n15062), .A2(n16044), .B1(n14634), .B2(n15060), .ZN(
        n3529) );
  OAI22_X1 U1487 ( .A1(n15062), .A2(n16043), .B1(n14640), .B2(n15060), .ZN(
        n3528) );
  OAI22_X1 U1488 ( .A1(n15086), .A2(n16033), .B1(n14714), .B2(n15079), .ZN(
        n3392) );
  OAI22_X1 U1489 ( .A1(n15082), .A2(n16030), .B1(n14633), .B2(n15079), .ZN(
        n3414) );
  OAI22_X1 U1490 ( .A1(n15087), .A2(n15932), .B1(n14660), .B2(n15079), .ZN(
        n1775) );
  OAI22_X1 U1491 ( .A1(n15105), .A2(n15922), .B1(n14659), .B2(n15100), .ZN(
        n1263) );
  OAI22_X1 U1492 ( .A1(n15190), .A2(n15745), .B1(n14654), .B2(n1085), .ZN(
        n1933) );
  OAI22_X1 U1493 ( .A1(n15012), .A2(n15638), .B1(n14681), .B2(n1119), .ZN(
        n1814) );
  OAI22_X1 U1494 ( .A1(n15008), .A2(n15630), .B1(n14621), .B2(n15000), .ZN(
        n1602) );
  OAI22_X1 U1495 ( .A1(n15002), .A2(n15624), .B1(n14705), .B2(n15001), .ZN(
        n1630) );
  OAI22_X1 U1496 ( .A1(n15212), .A2(n15614), .B1(n15220), .B2(n14620), .ZN(
        n1378) );
  OAI22_X1 U1497 ( .A1(n15212), .A2(n15610), .B1(n15218), .B2(n14686), .ZN(
        n1400) );
  OAI22_X1 U1498 ( .A1(n15006), .A2(n15597), .B1(n14645), .B2(n15000), .ZN(
        n1610) );
  OAI22_X1 U1499 ( .A1(n15014), .A2(n15566), .B1(n14669), .B2(n1119), .ZN(
        n1810) );
  OAI22_X1 U1500 ( .A1(n15067), .A2(n16116), .B1(n14636), .B2(n15060), .ZN(
        n1863) );
  OAI22_X1 U1501 ( .A1(n15107), .A2(n16082), .B1(n14631), .B2(n15099), .ZN(
        n1253) );
  OAI22_X1 U1502 ( .A1(n15103), .A2(n16079), .B1(n14677), .B2(n15099), .ZN(
        n3569) );
  OAI22_X1 U1503 ( .A1(n15063), .A2(n16040), .B1(n14664), .B2(n15060), .ZN(
        n3522) );
  OAI22_X1 U1504 ( .A1(n15064), .A2(n16036), .B1(n14668), .B2(n15060), .ZN(
        n3520) );
  OAI22_X1 U1505 ( .A1(n15082), .A2(n15952), .B1(n14641), .B2(n15079), .ZN(
        n3411) );
  OAI22_X1 U1506 ( .A1(n15104), .A2(n15933), .B1(n14713), .B2(n15100), .ZN(
        n3563) );
  OAI22_X1 U1507 ( .A1(n14976), .A2(n15767), .B1(n14631), .B2(n1124), .ZN(
        n1509) );
  OAI22_X1 U1508 ( .A1(n14973), .A2(n15764), .B1(n14667), .B2(n14968), .ZN(
        n1521) );
  OAI22_X1 U1509 ( .A1(n14972), .A2(n15763), .B1(n14679), .B2(n1124), .ZN(
        n1525) );
  OAI22_X1 U1510 ( .A1(n14971), .A2(n15762), .B1(n14697), .B2(n1124), .ZN(
        n1531) );
  OAI22_X1 U1511 ( .A1(n14969), .A2(n15755), .B1(n14712), .B2(n1124), .ZN(
        n1536) );
  OAI22_X1 U1512 ( .A1(n14973), .A2(n15754), .B1(n14715), .B2(n1124), .ZN(
        n1537) );
  OAI22_X1 U1513 ( .A1(n15007), .A2(n15753), .B1(n14630), .B2(n15000), .ZN(
        n1605) );
  OAI22_X1 U1514 ( .A1(n15191), .A2(n15737), .B1(n14633), .B2(n1085), .ZN(
        n1926) );
  OAI22_X1 U1515 ( .A1(n15191), .A2(n15736), .B1(n14639), .B2(n15184), .ZN(
        n1928) );
  OAI22_X1 U1516 ( .A1(n15188), .A2(n15735), .B1(n14672), .B2(n1085), .ZN(
        n1939) );
  OAI22_X1 U1517 ( .A1(n15211), .A2(n15685), .B1(n15220), .B2(n14629), .ZN(
        n1381) );
  OAI22_X1 U1518 ( .A1(n15007), .A2(n15629), .B1(n14636), .B2(n15000), .ZN(
        n1607) );
  OAI22_X1 U1519 ( .A1(n15004), .A2(n15627), .B1(n14675), .B2(n15001), .ZN(
        n1620) );
  OAI22_X1 U1520 ( .A1(n15003), .A2(n15626), .B1(n14687), .B2(n15001), .ZN(
        n1624) );
  OAI22_X1 U1521 ( .A1(n15003), .A2(n15625), .B1(n14693), .B2(n15000), .ZN(
        n1626) );
  OAI22_X1 U1522 ( .A1(n15211), .A2(n15612), .B1(n15219), .B2(n14635), .ZN(
        n1383) );
  OAI22_X1 U1523 ( .A1(n15212), .A2(n15609), .B1(n15218), .B2(n14692), .ZN(
        n1402) );
  OAI22_X1 U1524 ( .A1(n15212), .A2(n15608), .B1(n15217), .B2(n14704), .ZN(
        n1406) );
  OAI22_X1 U1525 ( .A1(n15012), .A2(n15565), .B1(n14690), .B2(n1119), .ZN(
        n1817) );
  OAI22_X1 U1526 ( .A1(n15002), .A2(n15559), .B1(n14708), .B2(n15001), .ZN(
        n1631) );
  OAI22_X1 U1527 ( .A1(n15187), .A2(n15552), .B1(n14689), .B2(n1085), .ZN(
        n3774) );
  OAI22_X1 U1528 ( .A1(n15006), .A2(n15543), .B1(n14642), .B2(n15000), .ZN(
        n1609) );
  OAI22_X1 U1529 ( .A1(n15185), .A2(n15456), .B1(n14680), .B2(n1085), .ZN(
        n3775) );
  OAI22_X1 U1530 ( .A1(n15010), .A2(n15534), .B1(n14711), .B2(n1119), .ZN(
        n1824) );
  OAI22_X1 U1531 ( .A1(n15103), .A2(n16078), .B1(n14695), .B2(n15100), .ZN(
        n3568) );
  OAI22_X1 U1532 ( .A1(n15104), .A2(n15934), .B1(n14710), .B2(n15100), .ZN(
        n3564) );
  OAI22_X1 U1533 ( .A1(n15016), .A2(n15673), .B1(n14642), .B2(n15009), .ZN(
        n1801) );
  OAI22_X1 U1534 ( .A1(n15015), .A2(n15672), .B1(n14645), .B2(n15009), .ZN(
        n1802) );
  OAI22_X1 U1535 ( .A1(n15015), .A2(n15671), .B1(n14648), .B2(n1119), .ZN(
        n1803) );
  OAI22_X1 U1536 ( .A1(n15192), .A2(n15637), .B1(n1085), .B2(n14626), .ZN(
        n1924) );
  OAI22_X1 U1537 ( .A1(n15190), .A2(n15636), .B1(n1085), .B2(n14650), .ZN(
        n1932) );
  OAI22_X1 U1538 ( .A1(n15187), .A2(n15635), .B1(n1085), .B2(n14698), .ZN(
        n1948) );
  OAI22_X1 U1539 ( .A1(n15186), .A2(n15634), .B1(n1085), .B2(n14701), .ZN(
        n1949) );
  OAI22_X1 U1540 ( .A1(n15212), .A2(n15633), .B1(n15219), .B2(n14659), .ZN(
        n1391) );
  OAI22_X1 U1541 ( .A1(n15017), .A2(n15623), .B1(n14627), .B2(n1119), .ZN(
        n1796) );
  OAI22_X1 U1542 ( .A1(n15015), .A2(n15622), .B1(n14651), .B2(n1119), .ZN(
        n1804) );
  OAI22_X1 U1543 ( .A1(n15011), .A2(n15621), .B1(n14699), .B2(n15009), .ZN(
        n1820) );
  OAI22_X1 U1544 ( .A1(n15011), .A2(n15620), .B1(n14702), .B2(n1119), .ZN(
        n1821) );
  OAI22_X1 U1545 ( .A1(n15191), .A2(n15619), .B1(n14642), .B2(n1085), .ZN(
        n1929) );
  OAI22_X1 U1546 ( .A1(n15190), .A2(n15618), .B1(n14645), .B2(n1085), .ZN(
        n1930) );
  OAI22_X1 U1547 ( .A1(n15189), .A2(n15617), .B1(n1085), .B2(n14665), .ZN(
        n1937) );
  OAI22_X1 U1548 ( .A1(n15189), .A2(n15615), .B1(n1085), .B2(n14695), .ZN(
        n1947) );
  OAI22_X1 U1549 ( .A1(n15017), .A2(n15596), .B1(n14621), .B2(n1119), .ZN(
        n1794) );
  OAI22_X1 U1550 ( .A1(n15016), .A2(n15595), .B1(n14633), .B2(n15009), .ZN(
        n1798) );
  OAI22_X1 U1551 ( .A1(n15016), .A2(n15594), .B1(n14636), .B2(n1119), .ZN(
        n1799) );
  OAI22_X1 U1552 ( .A1(n15016), .A2(n15593), .B1(n14639), .B2(n15009), .ZN(
        n1800) );
  OAI22_X1 U1553 ( .A1(n15013), .A2(n15592), .B1(n14672), .B2(n1119), .ZN(
        n1811) );
  OAI22_X1 U1554 ( .A1(n15011), .A2(n15588), .B1(n14705), .B2(n1119), .ZN(
        n1822) );
  OAI22_X1 U1555 ( .A1(n15011), .A2(n15564), .B1(n14708), .B2(n1119), .ZN(
        n1823) );
  OAI22_X1 U1556 ( .A1(n15190), .A2(n15563), .B1(n14648), .B2(n1085), .ZN(
        n1931) );
  OAI22_X1 U1557 ( .A1(n15191), .A2(n15556), .B1(n1085), .B2(n14635), .ZN(
        n1927) );
  OAI22_X1 U1558 ( .A1(n15188), .A2(n15554), .B1(n15184), .B2(n14674), .ZN(
        n1940) );
  OAI22_X1 U1559 ( .A1(n15187), .A2(n15553), .B1(n15184), .B2(n14686), .ZN(
        n1944) );
  OAI22_X1 U1560 ( .A1(n15187), .A2(n15551), .B1(n15184), .B2(n14692), .ZN(
        n1946) );
  OAI22_X1 U1561 ( .A1(n15186), .A2(n15550), .B1(n1085), .B2(n14704), .ZN(
        n1950) );
  OAI22_X1 U1562 ( .A1(n15014), .A2(n15533), .B1(n14714), .B2(n1119), .ZN(
        n1825) );
  OAI22_X1 U1563 ( .A1(n15212), .A2(n15440), .B1(n15216), .B2(n14710), .ZN(
        n1408) );
  OAI22_X1 U1564 ( .A1(n15212), .A2(n15439), .B1(n15216), .B2(n14713), .ZN(
        n1409) );
  OAI22_X1 U1565 ( .A1(n15185), .A2(n15431), .B1(n1085), .B2(n14710), .ZN(
        n3729) );
  OAI22_X1 U1566 ( .A1(n15186), .A2(n15430), .B1(n1085), .B2(n14713), .ZN(
        n3728) );
  OAI22_X1 U1567 ( .A1(n15068), .A2(n16119), .B1(n14621), .B2(n15060), .ZN(
        n1858) );
  OAI22_X1 U1568 ( .A1(n15063), .A2(n16041), .B1(n14660), .B2(n15060), .ZN(
        n3523) );
  OAI22_X1 U1569 ( .A1(n15064), .A2(n16035), .B1(n14690), .B2(n15061), .ZN(
        n3517) );
  OAI22_X1 U1570 ( .A1(n15082), .A2(n15951), .B1(n14644), .B2(n15079), .ZN(
        n3410) );
  OAI22_X1 U1571 ( .A1(n15188), .A2(n15616), .B1(n15184), .B2(n14677), .ZN(
        n1941) );
  OAI22_X1 U1572 ( .A1(n15212), .A2(n15613), .B1(n15220), .B2(n14624), .ZN(
        n1379) );
  OAI22_X1 U1573 ( .A1(n15013), .A2(n15591), .B1(n14675), .B2(n1119), .ZN(
        n1812) );
  OAI22_X1 U1574 ( .A1(n15013), .A2(n15590), .B1(n14687), .B2(n1119), .ZN(
        n1816) );
  OAI22_X1 U1575 ( .A1(n15012), .A2(n15589), .B1(n14693), .B2(n1119), .ZN(
        n1818) );
  OAI22_X1 U1576 ( .A1(n15189), .A2(n15587), .B1(n15184), .B2(n14659), .ZN(
        n3777) );
  OAI22_X1 U1577 ( .A1(n15192), .A2(n15557), .B1(n1085), .B2(n14620), .ZN(
        n1922) );
  OAI22_X1 U1578 ( .A1(n15017), .A2(n15535), .B1(n14630), .B2(n15009), .ZN(
        n1797) );
  OAI22_X1 U1579 ( .A1(n15192), .A2(n15532), .B1(n1085), .B2(n14623), .ZN(
        n1923) );
  OAI22_X1 U1580 ( .A1(n15192), .A2(n15508), .B1(n1085), .B2(n14629), .ZN(
        n1925) );
  OAI22_X1 U1581 ( .A1(n15211), .A2(n15444), .B1(n15220), .B2(n14626), .ZN(
        n1380) );
  OAI22_X1 U1582 ( .A1(n15212), .A2(n15443), .B1(n15219), .B2(n14650), .ZN(
        n1388) );
  OAI22_X1 U1583 ( .A1(n15212), .A2(n15442), .B1(n15217), .B2(n14698), .ZN(
        n1404) );
  OAI22_X1 U1584 ( .A1(n15212), .A2(n15441), .B1(n15217), .B2(n14701), .ZN(
        n1405) );
  NOR3_X1 U1585 ( .A1(n15304), .A2(Write_address[1]), .A3(n15312), .ZN(n1109)
         );
  NOR3_X1 U1586 ( .A1(n15304), .A2(Write_address[2]), .A3(n15311), .ZN(n1113)
         );
  NOR3_X1 U1587 ( .A1(Write_address[1]), .A2(Write_address[2]), .A3(
        Write_address[0]), .ZN(n1117) );
  NOR3_X1 U1588 ( .A1(Write_address[0]), .A2(Write_address[2]), .A3(n15311), 
        .ZN(n1114) );
  NOR3_X1 U1589 ( .A1(n15311), .A2(Write_address[0]), .A3(n15312), .ZN(n1108)
         );
  NOR3_X1 U1590 ( .A1(Write_address[1]), .A2(Write_address[2]), .A3(n15304), 
        .ZN(n1115) );
  NOR3_X1 U1591 ( .A1(Write_address[0]), .A2(Write_address[1]), .A3(n15312), 
        .ZN(n1111) );
  AOI21_X1 U1592 ( .B1(n1117), .B2(n3056), .A(n16314), .ZN(n2580) );
  NOR2_X1 U1593 ( .A1(Write_address[3]), .A2(Write_address[4]), .ZN(n3056) );
  INV_X1 U1594 ( .A(Write_address[1]), .ZN(n15311) );
  INV_X1 U1595 ( .A(Write_address[2]), .ZN(n15312) );
  INV_X1 U1596 ( .A(Write_address[0]), .ZN(n15304) );
  AND4_X1 U1597 ( .A1(n3048), .A2(n2580), .A3(n3049), .A4(n3050), .ZN(n1167)
         );
  NOR3_X1 U1598 ( .A1(n3051), .A2(n3052), .A3(n3054), .ZN(n3050) );
  INV_X1 U1599 ( .A(Data_in[0]), .ZN(n15315) );
  INV_X1 U1600 ( .A(Data_in[5]), .ZN(n15320) );
  INV_X1 U1601 ( .A(Data_in[18]), .ZN(n15333) );
  INV_X1 U1602 ( .A(Data_in[22]), .ZN(n15337) );
  INV_X1 U1603 ( .A(Data_in[24]), .ZN(n15339) );
  INV_X1 U1604 ( .A(Data_in[28]), .ZN(n15343) );
  INV_X1 U1605 ( .A(Data_in[14]), .ZN(n15329) );
  INV_X1 U1606 ( .A(Data_in[13]), .ZN(n15328) );
  INV_X1 U1607 ( .A(Data_in[9]), .ZN(n15324) );
  INV_X1 U1608 ( .A(Data_in[4]), .ZN(n15319) );
  INV_X1 U1609 ( .A(Data_in[6]), .ZN(n15321) );
  INV_X1 U1610 ( .A(Data_in[17]), .ZN(n15332) );
  INV_X1 U1611 ( .A(Data_in[20]), .ZN(n15335) );
  INV_X1 U1612 ( .A(Data_in[11]), .ZN(n15326) );
  INV_X1 U1613 ( .A(Data_in[12]), .ZN(n15327) );
  INV_X1 U1614 ( .A(Data_in[21]), .ZN(n15336) );
  INV_X1 U1615 ( .A(Data_in[29]), .ZN(n15344) );
  INV_X1 U1616 ( .A(Data_in[16]), .ZN(n15331) );
  INV_X1 U1617 ( .A(Data_in[19]), .ZN(n15334) );
  INV_X1 U1618 ( .A(Data_in[2]), .ZN(n15317) );
  INV_X1 U1619 ( .A(Data_in[3]), .ZN(n15318) );
  INV_X1 U1620 ( .A(Data_in[1]), .ZN(n15316) );
  INV_X1 U1621 ( .A(Data_in[7]), .ZN(n15322) );
  INV_X1 U1622 ( .A(Data_in[8]), .ZN(n15323) );
  INV_X1 U1623 ( .A(Data_in[10]), .ZN(n15325) );
  INV_X1 U1624 ( .A(Data_in[15]), .ZN(n15330) );
  INV_X1 U1625 ( .A(Data_in[23]), .ZN(n15338) );
  INV_X1 U1626 ( .A(Data_in[25]), .ZN(n15340) );
  INV_X1 U1627 ( .A(Data_in[26]), .ZN(n15341) );
  INV_X1 U1628 ( .A(Data_in[27]), .ZN(n15342) );
  INV_X1 U1629 ( .A(Data_in[30]), .ZN(n15345) );
  INV_X1 U1630 ( .A(Data_in[31]), .ZN(n15346) );
  INV_X1 U1631 ( .A(Write_address[3]), .ZN(n15313) );
  INV_X1 U1632 ( .A(Write_address[4]), .ZN(n15314) );
  NOR3_X1 U1633 ( .A1(n2583), .A2(n2584), .A3(n2585), .ZN(n2582) );
  OAI22_X1 U1634 ( .A1(n9389), .A2(n14750), .B1(n9768), .B2(n14760), .ZN(n2262) );
  OAI21_X1 U1635 ( .B1(n9664), .B2(n1471), .A(n15275), .ZN(n2263) );
  OAI22_X1 U1636 ( .A1(n9827), .A2(n14829), .B1(n9417), .B2(n14785), .ZN(n2260) );
  OAI22_X1 U1637 ( .A1(n9400), .A2(n14762), .B1(n3909), .B2(n14752), .ZN(n2317) );
  OAI211_X1 U1638 ( .C1(n14763), .C2(n15463), .A(n15272), .B(n2319), .ZN(n2312) );
  OAI222_X1 U1639 ( .A1(n3256), .A2(n14793), .B1(n9563), .B2(n14816), .C1(
        n3956), .C2(n1471), .ZN(n2314) );
  OAI22_X1 U1640 ( .A1(n3869), .A2(n14829), .B1(n3323), .B2(n14785), .ZN(n1712) );
  OAI22_X1 U1641 ( .A1(n3143), .A2(n14829), .B1(n3973), .B2(n1634), .ZN(n1718)
         );
  OAI21_X1 U1642 ( .B1(n3837), .B2(n14811), .A(n1720), .ZN(n1716) );
  OAI22_X1 U1643 ( .A1(n3645), .A2(n14829), .B1(n3322), .B2(n14785), .ZN(n1449) );
  OAI22_X1 U1644 ( .A1(n3144), .A2(n14829), .B1(n3974), .B2(n1634), .ZN(n1463)
         );
  OAI21_X1 U1645 ( .B1(n3815), .B2(n14811), .A(n1647), .ZN(n1454) );
  OAI22_X1 U1646 ( .A1(n14788), .A2(n15388), .B1(n3243), .B2(n14796), .ZN(
        n2243) );
  OAI221_X1 U1647 ( .B1(n9821), .B2(n1471), .C1(n9843), .C2(n14753), .A(n2248), 
        .ZN(n2241) );
  OAI22_X1 U1648 ( .A1(n3084), .A2(n14811), .B1(n9771), .B2(n14717), .ZN(n2246) );
  OAI22_X1 U1649 ( .A1(n14788), .A2(n15384), .B1(n3258), .B2(n14796), .ZN(
        n2106) );
  OAI221_X1 U1650 ( .B1(n9823), .B2(n1471), .C1(n9844), .C2(n14754), .A(n2111), 
        .ZN(n2104) );
  OAI22_X1 U1651 ( .A1(n3707), .A2(n14811), .B1(n9773), .B2(n14717), .ZN(n2109) );
  OAI22_X1 U1652 ( .A1(n14789), .A2(n15385), .B1(n3244), .B2(n14796), .ZN(
        n2167) );
  OAI221_X1 U1653 ( .B1(n9822), .B2(n1471), .C1(n9845), .C2(n14754), .A(n2172), 
        .ZN(n2165) );
  OAI22_X1 U1654 ( .A1(n3085), .A2(n14811), .B1(n9772), .B2(n14717), .ZN(n2170) );
  OAI22_X1 U1655 ( .A1(n14788), .A2(n15391), .B1(n3239), .B2(n14795), .ZN(
        n2478) );
  OAI221_X1 U1656 ( .B1(n9819), .B2(n14828), .C1(n9842), .C2(n14753), .A(n2483), .ZN(n2476) );
  OAI22_X1 U1657 ( .A1(n3079), .A2(n14811), .B1(n9770), .B2(n14717), .ZN(n2481) );
  OAI22_X1 U1658 ( .A1(n14789), .A2(n15392), .B1(n3236), .B2(n14795), .ZN(
        n2570) );
  OAI221_X1 U1659 ( .B1(n9816), .B2(n1471), .C1(n9841), .C2(n14753), .A(n2575), 
        .ZN(n2568) );
  OAI22_X1 U1660 ( .A1(n3708), .A2(n14811), .B1(n9769), .B2(n14717), .ZN(n2573) );
  OAI22_X1 U1661 ( .A1(n14789), .A2(n15383), .B1(n3245), .B2(n14795), .ZN(
        n1845) );
  OAI221_X1 U1662 ( .B1(n9824), .B2(n1471), .C1(n9846), .C2(n14754), .A(n1852), 
        .ZN(n1843) );
  OAI22_X1 U1663 ( .A1(n3706), .A2(n14811), .B1(n9774), .B2(n14717), .ZN(n1850) );
  AOI222_X1 U1664 ( .A1(n1771), .A2(n3070), .B1(n1772), .B2(n1773), .C1(n15293), .C2(n1774), .ZN(n1770) );
  AOI221_X1 U1665 ( .B1(n14719), .B2(n16124), .C1(n14808), .C2(n16269), .A(
        n1786), .ZN(n1773) );
  AOI211_X1 U1666 ( .C1(n14819), .C2(n15510), .A(n1787), .B(n1788), .ZN(n1772)
         );
  OAI222_X1 U1667 ( .A1(n16068), .A2(n1835), .B1(n15898), .B2(n1836), .C1(
        n3375), .C2(n1839), .ZN(n2308) );
  OAI222_X1 U1668 ( .A1(n16071), .A2(n1835), .B1(n15903), .B2(n1836), .C1(
        n3372), .C2(n1839), .ZN(n2490) );
  OAI222_X1 U1669 ( .A1(n16145), .A2(n1835), .B1(n15897), .B2(n1836), .C1(
        n3379), .C2(n1839), .ZN(n2255) );
  OAI222_X1 U1670 ( .A1(n16070), .A2(n1835), .B1(n15901), .B2(n1836), .C1(
        n3373), .C2(n1839), .ZN(n2455) );
  AOI222_X1 U1671 ( .A1(n3929), .A2(n14737), .B1(n9341), .B2(n14803), .C1(
        n14746), .C2(n15854), .ZN(n2319) );
  AOI222_X1 U1672 ( .A1(n3242), .A2(n14747), .B1(n14842), .B2(n15729), .C1(
        n14741), .C2(n16151), .ZN(n2334) );
  OAI222_X1 U1673 ( .A1(n9334), .A2(n14756), .B1(n3343), .B2(n14816), .C1(
        n9364), .C2(n14763), .ZN(n1763) );
  AOI221_X1 U1674 ( .B1(n14835), .B2(n16044), .C1(n14740), .C2(n15578), .A(
        n2500), .ZN(n2494) );
  OAI222_X1 U1675 ( .A1(n9478), .A2(n14799), .B1(n3861), .B2(n14816), .C1(
        n9396), .C2(n14763), .ZN(n2500) );
  OAI222_X1 U1676 ( .A1(n3839), .A2(n14828), .B1(n3720), .B2(n14732), .C1(
        n14795), .C2(n15488), .ZN(n2282) );
  OAI222_X1 U1677 ( .A1(n3855), .A2(n14828), .B1(n3718), .B2(n14732), .C1(
        n14795), .C2(n15485), .ZN(n2152) );
  OAI222_X1 U1678 ( .A1(n3269), .A2(n14793), .B1(n3703), .B2(n14732), .C1(
        n3961), .C2(n14763), .ZN(n2211) );
  AOI211_X1 U1679 ( .C1(n14723), .C2(n15980), .A(n2530), .B(n15270), .ZN(n2527) );
  OAI222_X1 U1680 ( .A1(n3685), .A2(n14816), .B1(n9659), .B2(n14732), .C1(
        n3213), .C2(n14792), .ZN(n2530) );
  AOI211_X1 U1681 ( .C1(n14723), .C2(n15977), .A(n2385), .B(n15270), .ZN(n2382) );
  OAI222_X1 U1682 ( .A1(n3951), .A2(n14815), .B1(n9660), .B2(n14732), .C1(
        n3214), .C2(n14792), .ZN(n2385) );
  AOI211_X1 U1683 ( .C1(n14722), .C2(n15975), .A(n1965), .B(n15269), .ZN(n1953) );
  OAI222_X1 U1684 ( .A1(n3921), .A2(n14814), .B1(n9661), .B2(n14732), .C1(
        n3215), .C2(n14793), .ZN(n1965) );
  AOI211_X1 U1685 ( .C1(n14722), .C2(n15974), .A(n1871), .B(n15270), .ZN(n1866) );
  OAI222_X1 U1686 ( .A1(n3922), .A2(n14814), .B1(n9662), .B2(n14732), .C1(
        n3230), .C2(n14792), .ZN(n1871) );
  OAI222_X1 U1687 ( .A1(n2328), .A2(n2329), .B1(n2330), .B2(n2331), .C1(n2332), 
        .C2(n2333), .ZN(n2327) );
  OAI221_X1 U1688 ( .B1(n9562), .B2(n14755), .C1(n9854), .C2(n1471), .A(n2339), 
        .ZN(n2328) );
  OAI221_X1 U1689 ( .B1(n3267), .B2(n14790), .C1(n3917), .C2(n14761), .A(n2335), .ZN(n2332) );
  OAI211_X1 U1690 ( .C1(n14799), .C2(n15492), .A(n15271), .B(n2334), .ZN(n2333) );
  AOI221_X1 U1691 ( .B1(n2180), .B2(n2344), .C1(n2345), .C2(n2346), .A(n2347), 
        .ZN(n2343) );
  AOI221_X1 U1692 ( .B1(n14721), .B2(n16126), .C1(n9722), .C2(n14832), .A(
        n2352), .ZN(n2346) );
  AOI211_X1 U1693 ( .C1(n3931), .C2(n14802), .A(n2353), .B(n2354), .ZN(n2345)
         );
  AOI21_X1 U1694 ( .B1(n2348), .B2(n2349), .A(n2187), .ZN(n2347) );
  AOI221_X1 U1695 ( .B1(n2180), .B2(n2363), .C1(n2364), .C2(n2365), .A(n2366), 
        .ZN(n2362) );
  AOI221_X1 U1696 ( .B1(n14721), .B2(n16127), .C1(n9721), .C2(n14832), .A(
        n2371), .ZN(n2365) );
  AOI211_X1 U1697 ( .C1(n3930), .C2(n14802), .A(n2372), .B(n2373), .ZN(n2364)
         );
  AOI21_X1 U1698 ( .B1(n2367), .B2(n2368), .A(n2187), .ZN(n2366) );
  AOI221_X1 U1699 ( .B1(n2180), .B2(n2181), .C1(n2182), .C2(n2183), .A(n2184), 
        .ZN(n2179) );
  AOI221_X1 U1700 ( .B1(n14719), .B2(n16125), .C1(n9723), .C2(n14830), .A(
        n2190), .ZN(n2183) );
  AOI211_X1 U1701 ( .C1(n3932), .C2(n14801), .A(n2191), .B(n2192), .ZN(n2182)
         );
  AOI21_X1 U1702 ( .B1(n2185), .B2(n2186), .A(n2187), .ZN(n2184) );
  AOI221_X1 U1703 ( .B1(n14818), .B2(n15581), .C1(n14725), .C2(n16037), .A(
        Read_one_address[1]), .ZN(n2335) );
  OAI222_X1 U1704 ( .A1(n3340), .A2(n14814), .B1(n9775), .B2(n1670), .C1(n9388), .C2(n14798), .ZN(n1777) );
  OAI222_X1 U1705 ( .A1(n3119), .A2(n14815), .B1(n9785), .B2(n14718), .C1(
        n9652), .C2(n14731), .ZN(n2242) );
  OAI222_X1 U1706 ( .A1(n3121), .A2(n14814), .B1(n9787), .B2(n1670), .C1(n9651), .C2(n14731), .ZN(n2105) );
  OAI222_X1 U1707 ( .A1(n3120), .A2(n14815), .B1(n9786), .B2(n14718), .C1(
        n9648), .C2(n14731), .ZN(n2166) );
  OAI222_X1 U1708 ( .A1(n3118), .A2(n14816), .B1(n9784), .B2(n14718), .C1(
        n9653), .C2(n14731), .ZN(n2477) );
  OAI222_X1 U1709 ( .A1(n3968), .A2(n14763), .B1(n14752), .B2(n15461), .C1(
        n3324), .C2(n14731), .ZN(n1704) );
  OAI222_X1 U1710 ( .A1(n3969), .A2(n14763), .B1(n14752), .B2(n15460), .C1(
        n3325), .C2(n14731), .ZN(n1441) );
  OAI222_X1 U1711 ( .A1(n14762), .A2(n15358), .B1(n9384), .B2(n14797), .C1(
        n3889), .C2(n14731), .ZN(n2245) );
  OAI222_X1 U1712 ( .A1(n14762), .A2(n15356), .B1(n9386), .B2(n14799), .C1(
        n3919), .C2(n14731), .ZN(n2108) );
  OAI222_X1 U1713 ( .A1(n14762), .A2(n15357), .B1(n9385), .B2(n14799), .C1(
        n3899), .C2(n14731), .ZN(n2169) );
  OAI222_X1 U1714 ( .A1(n14762), .A2(n15359), .B1(n9383), .B2(n14799), .C1(
        n3818), .C2(n14731), .ZN(n2480) );
  OAI222_X1 U1715 ( .A1(n14762), .A2(n15361), .B1(n9382), .B2(n14797), .C1(
        n3666), .C2(n14731), .ZN(n2572) );
  OAI222_X1 U1716 ( .A1(n14762), .A2(n15355), .B1(n9387), .B2(n14797), .C1(
        n3925), .C2(n14731), .ZN(n1849) );
  OAI222_X1 U1717 ( .A1(n3826), .A2(n14815), .B1(n9779), .B2(n14718), .C1(
        n9480), .C2(n14799), .ZN(n2316) );
  OAI222_X1 U1718 ( .A1(n3117), .A2(n14814), .B1(n9783), .B2(n14718), .C1(
        n9650), .C2(n14732), .ZN(n2569) );
  OAI222_X1 U1719 ( .A1(n3122), .A2(n14814), .B1(n9788), .B2(n1670), .C1(n9649), .C2(n14732), .ZN(n1844) );
  AOI221_X1 U1720 ( .B1(n14747), .B2(n15826), .C1(n14770), .C2(n15877), .A(
        n2230), .ZN(n2229) );
  OAI222_X1 U1721 ( .A1(n3137), .A2(n14815), .B1(n9747), .B2(n14718), .C1(
        n3184), .C2(n14799), .ZN(n2230) );
  AOI221_X1 U1722 ( .B1(n14746), .B2(n15831), .C1(n14770), .C2(n15884), .A(
        n2519), .ZN(n2518) );
  OAI222_X1 U1723 ( .A1(n3858), .A2(n14815), .B1(n14717), .B2(n15464), .C1(
        n3139), .C2(n14799), .ZN(n2519) );
  AOI221_X1 U1724 ( .B1(n14747), .B2(n15829), .C1(n14769), .C2(n15882), .A(
        n2429), .ZN(n2428) );
  OAI222_X1 U1725 ( .A1(n3866), .A2(n14815), .B1(n14717), .B2(n15462), .C1(
        n3295), .C2(n14828), .ZN(n2429) );
  AOI221_X1 U1726 ( .B1(n14746), .B2(n15828), .C1(n14769), .C2(n15881), .A(
        n2392), .ZN(n2391) );
  OAI222_X1 U1727 ( .A1(n3671), .A2(n14815), .B1(n9751), .B2(n14718), .C1(
        n3821), .C2(n14799), .ZN(n2392) );
  AOI221_X1 U1728 ( .B1(n14747), .B2(n15827), .C1(n14769), .C2(n15880), .A(
        n2301), .ZN(n2300) );
  OAI222_X1 U1729 ( .A1(n3136), .A2(n14815), .B1(n9746), .B2(n14718), .C1(
        n3142), .C2(n14799), .ZN(n2301) );
  AOI221_X1 U1730 ( .B1(n14747), .B2(n15825), .C1(n14770), .C2(n15875), .A(
        n2089), .ZN(n2088) );
  OAI222_X1 U1731 ( .A1(n3669), .A2(n14814), .B1(n9749), .B2(n14718), .C1(
        n3185), .C2(n14798), .ZN(n2089) );
  AOI221_X1 U1732 ( .B1(n14746), .B2(n15824), .C1(n14771), .C2(n15874), .A(
        n2050), .ZN(n1982) );
  OAI222_X1 U1733 ( .A1(n3138), .A2(n14814), .B1(n9748), .B2(n1670), .C1(n3188), .C2(n14798), .ZN(n2050) );
  AOI221_X1 U1734 ( .B1(n14747), .B2(n15823), .C1(n14769), .C2(n15873), .A(
        n1885), .ZN(n1884) );
  OAI222_X1 U1735 ( .A1(n3667), .A2(n14814), .B1(n9750), .B2(n1670), .C1(n3189), .C2(n14798), .ZN(n1885) );
  AOI221_X1 U1736 ( .B1(n14734), .B2(n16238), .C1(n14748), .C2(n15820), .A(
        n2222), .ZN(n2221) );
  OAI221_X1 U1737 ( .B1(n3726), .B2(n1670), .C1(n3314), .C2(n14761), .A(n14844), .ZN(n2222) );
  AOI221_X1 U1738 ( .B1(n14835), .B2(n15623), .C1(n7821), .C2(n14747), .A(
        n2529), .ZN(n2528) );
  OAI221_X1 U1739 ( .B1(n9847), .B2(n14797), .C1(n9337), .C2(n14761), .A(
        n14844), .ZN(n2529) );
  AOI221_X1 U1740 ( .B1(n14834), .B2(n15622), .C1(n7822), .C2(n14746), .A(
        n2384), .ZN(n2383) );
  OAI221_X1 U1741 ( .B1(n9848), .B2(n14797), .C1(n9338), .C2(n14761), .A(
        n14844), .ZN(n2384) );
  AOI221_X1 U1742 ( .B1(n14735), .B2(n16239), .C1(n14748), .C2(n15821), .A(
        n2293), .ZN(n2292) );
  OAI221_X1 U1743 ( .B1(n3672), .B2(n14718), .C1(n3308), .C2(n14761), .A(
        n14844), .ZN(n2293) );
  AOI221_X1 U1744 ( .B1(n14833), .B2(n15621), .C1(n8085), .C2(n14746), .A(
        n1959), .ZN(n1954) );
  OAI221_X1 U1745 ( .B1(n9849), .B2(n14798), .C1(n9339), .C2(n14761), .A(
        n14844), .ZN(n1959) );
  AOI221_X1 U1746 ( .B1(n14834), .B2(n15620), .C1(n8086), .C2(n14746), .A(
        n1868), .ZN(n1867) );
  OAI221_X1 U1747 ( .B1(n9850), .B2(n14797), .C1(n9340), .C2(n14761), .A(
        n14844), .ZN(n1868) );
  AOI221_X1 U1748 ( .B1(n14747), .B2(n15832), .C1(n14770), .C2(n15885), .A(
        n2537), .ZN(n2536) );
  OAI222_X1 U1749 ( .A1(n3209), .A2(n14816), .B1(n9745), .B2(n1670), .C1(n3141), .C2(n14799), .ZN(n2537) );
  AOI221_X1 U1750 ( .B1(n14734), .B2(n16237), .C1(n14748), .C2(n15819), .A(
        n2078), .ZN(n2074) );
  OAI221_X1 U1751 ( .B1(n3796), .B2(n1670), .C1(n3316), .C2(n14760), .A(n14844), .ZN(n2078) );
  AOI221_X1 U1752 ( .B1(n14720), .B2(n9526), .C1(n14822), .C2(n15467), .A(
        n2369), .ZN(n2368) );
  OAI22_X1 U1753 ( .A1(n9447), .A2(n14750), .B1(n15993), .B2(n14796), .ZN(
        n2369) );
  AOI221_X1 U1754 ( .B1(n14720), .B2(n9523), .C1(n14822), .C2(n3091), .A(n2207), .ZN(n2206) );
  OAI22_X1 U1755 ( .A1(n15816), .A2(n14750), .B1(n15991), .B2(n14796), .ZN(
        n2207) );
  AOI221_X1 U1756 ( .B1(n14719), .B2(n9525), .C1(n14820), .C2(n15465), .A(
        n2188), .ZN(n2186) );
  OAI22_X1 U1757 ( .A1(n9446), .A2(n14749), .B1(n15990), .B2(n14796), .ZN(
        n2188) );
  AOI221_X1 U1758 ( .B1(n14747), .B2(n15769), .C1(n14768), .C2(n15847), .A(
        n2412), .ZN(n2407) );
  OAI222_X1 U1759 ( .A1(n3819), .A2(n14815), .B1(n9778), .B2(n1670), .C1(n9760), .C2(n14798), .ZN(n2412) );
  AOI221_X1 U1760 ( .B1(n14805), .B2(n16171), .C1(n14748), .C2(n15668), .A(
        n2558), .ZN(n2553) );
  OAI221_X1 U1761 ( .B1(n3807), .B2(n14718), .C1(n3962), .C2(n14811), .A(
        n15269), .ZN(n2558) );
  AOI221_X1 U1762 ( .B1(n14804), .B2(n16128), .C1(n14748), .C2(n15845), .A(
        n2410), .ZN(n2409) );
  OAI221_X1 U1763 ( .B1(n9811), .B2(n1670), .C1(n3094), .C2(n14812), .A(n15269), .ZN(n2410) );
  AOI221_X1 U1764 ( .B1(n14747), .B2(n15852), .C1(n9592), .C2(n14764), .A(
        n2556), .ZN(n2555) );
  OAI222_X1 U1765 ( .A1(n3854), .A2(n14816), .B1(n9500), .B2(n1670), .C1(n9472), .C2(n14799), .ZN(n2556) );
  AOI221_X1 U1766 ( .B1(n15291), .B2(n15417), .C1(n15292), .C2(n9604), .A(
        n1860), .ZN(n2354) );
  AOI221_X1 U1767 ( .B1(n15291), .B2(n15418), .C1(n15292), .C2(n9605), .A(
        n1860), .ZN(n2373) );
  AOI221_X1 U1768 ( .B1(n15291), .B2(n15413), .C1(n15292), .C2(n9606), .A(
        n1860), .ZN(n2192) );
  AOI211_X1 U1769 ( .C1(n3359), .C2(n14802), .A(n2250), .B(n2251), .ZN(n2238)
         );
  OAI21_X1 U1770 ( .B1(n3888), .B2(n14760), .A(n15274), .ZN(n2250) );
  AOI221_X1 U1771 ( .B1(n15291), .B2(n15414), .C1(n15292), .C2(n9598), .A(
        n1860), .ZN(n2251) );
  AOI211_X1 U1772 ( .C1(n3643), .C2(n14801), .A(n2113), .B(n2118), .ZN(n2099)
         );
  OAI21_X1 U1773 ( .B1(n3918), .B2(n14760), .A(n15273), .ZN(n2113) );
  AOI221_X1 U1774 ( .B1(n15291), .B2(n15410), .C1(n15292), .C2(n9599), .A(
        n1860), .ZN(n2118) );
  AOI211_X1 U1775 ( .C1(n3361), .C2(n14801), .A(n2174), .B(n2175), .ZN(n2162)
         );
  OAI21_X1 U1776 ( .B1(n3894), .B2(n14760), .A(n15275), .ZN(n2174) );
  AOI221_X1 U1777 ( .B1(n15291), .B2(n15412), .C1(n15292), .C2(n9600), .A(
        n1860), .ZN(n2175) );
  AOI211_X1 U1778 ( .C1(n14806), .C2(n16101), .A(n2268), .B(n2269), .ZN(n2256)
         );
  OAI21_X1 U1779 ( .B1(n3223), .B2(n14786), .A(n15275), .ZN(n2268) );
  AOI221_X1 U1780 ( .B1(n15291), .B2(n15415), .C1(n15292), .C2(n9608), .A(
        n1860), .ZN(n2269) );
  AOI211_X1 U1781 ( .C1(n3357), .C2(n14802), .A(n2485), .B(n2486), .ZN(n2473)
         );
  OAI21_X1 U1782 ( .B1(n3790), .B2(n14760), .A(n15276), .ZN(n2485) );
  AOI221_X1 U1783 ( .B1(n15291), .B2(n15422), .C1(n15292), .C2(n9601), .A(
        n1860), .ZN(n2486) );
  AOI211_X1 U1784 ( .C1(n3355), .C2(n14801), .A(n2577), .B(n2578), .ZN(n2565)
         );
  OAI21_X1 U1785 ( .B1(n3663), .B2(n14760), .A(n15276), .ZN(n2577) );
  AOI221_X1 U1786 ( .B1(n15291), .B2(n15425), .C1(n15292), .C2(n9602), .A(
        n1860), .ZN(n2578) );
  AOI211_X1 U1787 ( .C1(n3642), .C2(n14800), .A(n1856), .B(n1857), .ZN(n1840)
         );
  OAI21_X1 U1788 ( .B1(n3924), .B2(n14760), .A(n15273), .ZN(n1856) );
  AOI221_X1 U1789 ( .B1(n15291), .B2(n15407), .C1(n15292), .C2(n9603), .A(
        n1860), .ZN(n1857) );
  AOI221_X1 U1790 ( .B1(n14817), .B2(n15763), .C1(n9735), .C2(n14800), .A(
        n1873), .ZN(n2218) );
  AOI221_X1 U1791 ( .B1(n14818), .B2(n15764), .C1(n9734), .C2(n14800), .A(
        n1873), .ZN(n2289) );
  AOI221_X1 U1792 ( .B1(n14817), .B2(n15762), .C1(n9739), .C2(n14800), .A(
        n1873), .ZN(n2070) );
  AOI221_X1 U1793 ( .B1(n9434), .B2(n14748), .C1(n14771), .C2(n15698), .A(
        n1766), .ZN(n1726) );
  OAI22_X1 U1794 ( .A1(n9684), .A2(n14795), .B1(n9356), .B2(n14717), .ZN(n1766) );
  AOI221_X1 U1795 ( .B1(n9435), .B2(n14748), .C1(n14771), .C2(n15697), .A(
        n1697), .ZN(n1672) );
  OAI22_X1 U1796 ( .A1(n9685), .A2(n14795), .B1(n9357), .B2(n14717), .ZN(n1697) );
  AOI221_X1 U1797 ( .B1(n14782), .B2(n15662), .C1(n3225), .C2(n14831), .A(
        n2233), .ZN(n2226) );
  OAI22_X1 U1798 ( .A1(n3250), .A2(n14729), .B1(n9550), .B2(n14760), .ZN(n2233) );
  AOI221_X1 U1799 ( .B1(n14781), .B2(n15666), .C1(n3311), .C2(n14831), .A(
        n2540), .ZN(n2533) );
  OAI22_X1 U1800 ( .A1(n3247), .A2(n14729), .B1(n9548), .B2(n14760), .ZN(n2540) );
  AOI221_X1 U1801 ( .B1(n14781), .B2(n15665), .C1(n14842), .C2(n15840), .A(
        n2522), .ZN(n2515) );
  OAI22_X1 U1802 ( .A1(n3628), .A2(n14729), .B1(n9882), .B2(n14762), .ZN(n2522) );
  AOI221_X1 U1803 ( .B1(n14781), .B2(n15664), .C1(n3310), .C2(n14832), .A(
        n2395), .ZN(n2388) );
  OAI22_X1 U1804 ( .A1(n3248), .A2(n14730), .B1(n9552), .B2(n14759), .ZN(n2395) );
  AOI221_X1 U1805 ( .B1(n14782), .B2(n15663), .C1(n3203), .C2(n14832), .A(
        n2304), .ZN(n2297) );
  OAI22_X1 U1806 ( .A1(n3249), .A2(n14729), .B1(n9549), .B2(n14760), .ZN(n2304) );
  AOI221_X1 U1807 ( .B1(n14782), .B2(n15661), .C1(n3226), .C2(n14831), .A(
        n2092), .ZN(n2085) );
  OAI22_X1 U1808 ( .A1(n3251), .A2(n14729), .B1(n9553), .B2(n14759), .ZN(n2092) );
  AOI221_X1 U1809 ( .B1(n14781), .B2(n15660), .C1(n3227), .C2(n14831), .A(
        n2061), .ZN(n1975) );
  OAI22_X1 U1810 ( .A1(n3252), .A2(n14729), .B1(n9551), .B2(n14759), .ZN(n2061) );
  AOI221_X1 U1811 ( .B1(n14781), .B2(n15659), .C1(n3228), .C2(n14830), .A(
        n1935), .ZN(n1877) );
  OAI22_X1 U1812 ( .A1(n3253), .A2(n14729), .B1(n9554), .B2(n14759), .ZN(n1935) );
  AOI221_X1 U1813 ( .B1(n14737), .B2(n16086), .C1(n9448), .C2(n14746), .A(
        n2502), .ZN(n2492) );
  OAI221_X1 U1814 ( .B1(n3812), .B2(n14717), .C1(n3713), .C2(n14812), .A(
        n15269), .ZN(n2502) );
  AOI221_X1 U1815 ( .B1(n14736), .B2(n16085), .C1(n9449), .C2(n14746), .A(
        n2467), .ZN(n2457) );
  OAI221_X1 U1816 ( .B1(n3814), .B2(n1670), .C1(n3704), .C2(n14812), .A(n15269), .ZN(n2467) );
  AOI221_X1 U1817 ( .B1(n14781), .B2(n15667), .C1(n14841), .C2(n15841), .A(
        n2559), .ZN(n2552) );
  OAI22_X1 U1818 ( .A1(n3349), .A2(n14729), .B1(n9881), .B2(n14760), .ZN(n2559) );
  AOI221_X1 U1819 ( .B1(n14736), .B2(n15576), .C1(n14783), .C2(n15505), .A(
        n2413), .ZN(n2406) );
  OAI21_X1 U1820 ( .B1(n3296), .B2(n14828), .A(n2180), .ZN(n2413) );
  OAI221_X1 U1821 ( .B1(n9767), .B2(n14814), .C1(n3632), .C2(n14796), .A(n2450), .ZN(n2444) );
  AOI21_X1 U1822 ( .B1(n15300), .B2(n16009), .A(n2451), .ZN(n2450) );
  AOI221_X1 U1823 ( .B1(n3941), .B2(n1875), .C1(n3943), .C2(n14762), .A(n15298), .ZN(n2451) );
  OAI221_X1 U1824 ( .B1(n9766), .B2(n14813), .C1(n3633), .C2(n14796), .A(n2423), .ZN(n2417) );
  AOI21_X1 U1825 ( .B1(n15300), .B2(n16008), .A(n2424), .ZN(n2423) );
  AOI221_X1 U1826 ( .B1(n3946), .B2(n1875), .C1(n3947), .C2(n14760), .A(n15298), .ZN(n2424) );
  AOI221_X1 U1827 ( .B1(n14781), .B2(n15844), .C1(n3229), .C2(n14830), .A(
        n1765), .ZN(n1727) );
  OAI221_X1 U1828 ( .B1(n3148), .B2(n14813), .C1(n3873), .C2(n14730), .A(
        n15269), .ZN(n1765) );
  AOI221_X1 U1829 ( .B1(n14781), .B2(n15843), .C1(n3224), .C2(n14830), .A(
        n1696), .ZN(n1683) );
  OAI221_X1 U1830 ( .B1(n3149), .B2(n14813), .C1(n3649), .C2(n14730), .A(
        n15269), .ZN(n1696) );
  AOI221_X1 U1831 ( .B1(n15299), .B2(n15442), .C1(n14841), .C2(n15928), .A(
        n1966), .ZN(n1952) );
  OAI22_X1 U1832 ( .A1(n14797), .A2(n15351), .B1(n9614), .B2(n1652), .ZN(n1966) );
  AOI221_X1 U1833 ( .B1(n15299), .B2(n15441), .C1(n14842), .C2(n15927), .A(
        n1872), .ZN(n1865) );
  OAI22_X1 U1834 ( .A1(n14797), .A2(n15350), .B1(n9615), .B2(n1652), .ZN(n1872) );
  AOI221_X1 U1835 ( .B1(n14782), .B2(n15387), .C1(n14840), .C2(n9890), .A(
        n2208), .ZN(n2205) );
  OAI22_X1 U1836 ( .A1(n16216), .A2(n14729), .B1(n9506), .B2(n14760), .ZN(
        n2208) );
  AOI221_X1 U1837 ( .B1(n14781), .B2(n15386), .C1(n14841), .C2(n9869), .A(
        n2189), .ZN(n2185) );
  OAI22_X1 U1838 ( .A1(n16215), .A2(n14729), .B1(n3353), .B2(n14759), .ZN(
        n2189) );
  AOI221_X1 U1839 ( .B1(n14746), .B2(n15771), .C1(n14725), .C2(n15723), .A(
        n2501), .ZN(n2493) );
  OAI21_X1 U1840 ( .B1(n3132), .B2(n14786), .A(n2180), .ZN(n2501) );
  AOI221_X1 U1841 ( .B1(n14746), .B2(n15770), .C1(n14725), .C2(n15722), .A(
        n2466), .ZN(n2458) );
  OAI21_X1 U1842 ( .B1(n3133), .B2(n14787), .A(n2180), .ZN(n2466) );
  AOI211_X1 U1843 ( .C1(n14782), .C2(n15696), .A(n2503), .B(n2322), .ZN(n2491)
         );
  OAI222_X1 U1844 ( .A1(n3219), .A2(n14799), .B1(n9876), .B2(n14763), .C1(
        n9813), .C2(n1471), .ZN(n2503) );
  AOI211_X1 U1845 ( .C1(n14782), .C2(n15695), .A(n2468), .B(n2322), .ZN(n2456)
         );
  OAI222_X1 U1846 ( .A1(n3264), .A2(n14799), .B1(n9877), .B2(n14763), .C1(
        n9814), .C2(n14828), .ZN(n2468) );
  AOI211_X1 U1847 ( .C1(n14723), .C2(n16296), .A(n2321), .B(n2322), .ZN(n2309)
         );
  OAI222_X1 U1848 ( .A1(n3218), .A2(n14732), .B1(n3714), .B2(n14816), .C1(
        n3828), .C2(n14791), .ZN(n2321) );
  AOI211_X1 U1849 ( .C1(n3208), .C2(n14833), .A(n2411), .B(n2322), .ZN(n2408)
         );
  OAI222_X1 U1850 ( .A1(n3220), .A2(n14732), .B1(n9866), .B2(n14763), .C1(
        n3827), .C2(n14792), .ZN(n2411) );
  AOI211_X1 U1851 ( .C1(n14819), .C2(n15779), .A(n1873), .B(n2532), .ZN(n2525)
         );
  AOI221_X1 U1852 ( .B1(n3856), .B2(n1875), .C1(n3380), .C2(n14760), .A(n15298), .ZN(n2532) );
  AOI211_X1 U1853 ( .C1(n14819), .C2(n15778), .A(n1873), .B(n2387), .ZN(n2380)
         );
  AOI221_X1 U1854 ( .B1(n3820), .B2(n1875), .C1(n3664), .C2(n14760), .A(n15298), .ZN(n2387) );
  AOI211_X1 U1855 ( .C1(n14818), .C2(n15777), .A(n1873), .B(n1972), .ZN(n1945)
         );
  AOI221_X1 U1856 ( .B1(n3881), .B2(n1875), .C1(n3799), .C2(n14760), .A(n15298), .ZN(n1972) );
  AOI211_X1 U1857 ( .C1(n14818), .C2(n15776), .A(n1873), .B(n1874), .ZN(n1864)
         );
  AOI221_X1 U1858 ( .B1(n3884), .B2(n1875), .C1(n3801), .C2(n14760), .A(n15298), .ZN(n1874) );
  OAI221_X1 U1859 ( .B1(n9860), .B2(n14813), .C1(n14756), .C2(n15416), .A(
        n14618), .ZN(n2281) );
  OAI221_X1 U1860 ( .B1(n9861), .B2(n14814), .C1(n14757), .C2(n15411), .A(
        n14618), .ZN(n2151) );
  AOI221_X1 U1861 ( .B1(n14803), .B2(n16003), .C1(n3368), .C2(n14746), .A(
        n2232), .ZN(n2227) );
  OAI221_X1 U1862 ( .B1(n3830), .B2(n1670), .C1(n3174), .C2(n14813), .A(n15269), .ZN(n2232) );
  AOI221_X1 U1863 ( .B1(n14805), .B2(n16052), .C1(n14783), .C2(n15701), .A(
        n2431), .ZN(n2426) );
  OAI221_X1 U1864 ( .B1(n3201), .B2(n14716), .C1(n3150), .C2(n14812), .A(
        n15269), .ZN(n2431) );
  AOI221_X1 U1865 ( .B1(n14804), .B2(n16004), .C1(n3367), .C2(n14746), .A(
        n2303), .ZN(n2298) );
  OAI221_X1 U1866 ( .B1(n3829), .B2(n14718), .C1(n3171), .C2(n14813), .A(
        n15269), .ZN(n2303) );
  AOI221_X1 U1867 ( .B1(n14804), .B2(n16002), .C1(n3369), .C2(n14746), .A(
        n2091), .ZN(n2086) );
  OAI221_X1 U1868 ( .B1(n3834), .B2(n14717), .C1(n3177), .C2(n14813), .A(
        n15269), .ZN(n2091) );
  AOI221_X1 U1869 ( .B1(n14804), .B2(n16000), .C1(n3371), .C2(n14746), .A(
        n1889), .ZN(n1881) );
  OAI221_X1 U1870 ( .B1(n3836), .B2(n14717), .C1(n3192), .C2(n14812), .A(
        n15269), .ZN(n1889) );
  AOI221_X1 U1871 ( .B1(n14806), .B2(n16007), .C1(n3363), .C2(n14746), .A(
        n2539), .ZN(n2534) );
  OAI221_X1 U1872 ( .B1(n3809), .B2(n14718), .C1(n3125), .C2(n14813), .A(
        n15269), .ZN(n2539) );
  AOI221_X1 U1873 ( .B1(n14805), .B2(n16170), .C1(n3364), .C2(n14746), .A(
        n2521), .ZN(n2516) );
  OAI221_X1 U1874 ( .B1(n3810), .B2(n14718), .C1(n3126), .C2(n14812), .A(
        n15269), .ZN(n2521) );
  AOI221_X1 U1875 ( .B1(n14803), .B2(n16001), .C1(n3370), .C2(n14746), .A(
        n2059), .ZN(n1976) );
  OAI221_X1 U1876 ( .B1(n3835), .B2(n14718), .C1(n3187), .C2(n14812), .A(
        n15269), .ZN(n2059) );
  AOI221_X1 U1877 ( .B1(n14805), .B2(n16006), .C1(n3366), .C2(n14746), .A(
        n2394), .ZN(n2389) );
  OAI221_X1 U1878 ( .B1(n3207), .B2(n14717), .C1(n3168), .C2(n14812), .A(
        n15269), .ZN(n2394) );
  AOI221_X1 U1879 ( .B1(n14834), .B2(n15591), .C1(n14821), .C2(n15527), .A(
        n2249), .ZN(n2239) );
  OAI221_X1 U1880 ( .B1(n3233), .B2(n14790), .C1(n3156), .C2(n14718), .A(
        n14618), .ZN(n2249) );
  AOI221_X1 U1881 ( .B1(n14834), .B2(n15589), .C1(n14821), .C2(n15524), .A(
        n2112), .ZN(n2100) );
  OAI221_X1 U1882 ( .B1(n3235), .B2(n14791), .C1(n3159), .C2(n14718), .A(
        n14618), .ZN(n2112) );
  AOI221_X1 U1883 ( .B1(n14835), .B2(n15590), .C1(n14820), .C2(n15525), .A(
        n2173), .ZN(n2163) );
  OAI221_X1 U1884 ( .B1(n3234), .B2(n14791), .C1(n3158), .C2(n1670), .A(n14618), .ZN(n2173) );
  AOI221_X1 U1885 ( .B1(n14835), .B2(n15594), .C1(n14823), .C2(n15529), .A(
        n2484), .ZN(n2474) );
  OAI221_X1 U1886 ( .B1(n3232), .B2(n14790), .C1(n3153), .C2(n14718), .A(
        n14618), .ZN(n2484) );
  AOI221_X1 U1887 ( .B1(n14836), .B2(n15596), .C1(n14823), .C2(n15530), .A(
        n2576), .ZN(n2566) );
  OAI221_X1 U1888 ( .B1(n3712), .B2(n14791), .C1(n3711), .C2(n14717), .A(
        n14618), .ZN(n2576) );
  AOI221_X1 U1889 ( .B1(n14833), .B2(n15588), .C1(n14821), .C2(n15522), .A(
        n1854), .ZN(n1841) );
  OAI221_X1 U1890 ( .B1(n3710), .B2(n14790), .C1(n3709), .C2(n14717), .A(
        n14618), .ZN(n1854) );
  AOI211_X1 U1891 ( .C1(n14782), .C2(n16188), .A(n2082), .B(n15269), .ZN(n2072) );
  OAI222_X1 U1892 ( .A1(n3920), .A2(n14815), .B1(n3795), .B2(n14828), .C1(
        n9420), .C2(n14798), .ZN(n2082) );
  AOI211_X1 U1893 ( .C1(n14837), .C2(n16013), .A(n1764), .B(n15269), .ZN(n1737) );
  OAI22_X1 U1894 ( .A1(n9537), .A2(n14795), .B1(n9393), .B2(n14717), .ZN(n1764) );
  AOI211_X1 U1895 ( .C1(n14836), .C2(n16012), .A(n1694), .B(n15269), .ZN(n1684) );
  OAI22_X1 U1896 ( .A1(n9538), .A2(n14795), .B1(n9394), .B2(n14717), .ZN(n1694) );
  AOI211_X1 U1897 ( .C1(n14783), .C2(n16189), .A(n2223), .B(n15270), .ZN(n2220) );
  OAI222_X1 U1898 ( .A1(n3891), .A2(n14815), .B1(n3702), .B2(n14828), .C1(
        n9419), .C2(n14798), .ZN(n2223) );
  AOI211_X1 U1899 ( .C1(n14783), .C2(n16190), .A(n2294), .B(n15270), .ZN(n2291) );
  OAI222_X1 U1900 ( .A1(n3883), .A2(n14815), .B1(n3670), .B2(n1471), .C1(n9418), .C2(n14799), .ZN(n2294) );
  AOI211_X1 U1901 ( .C1(n9725), .C2(n14781), .A(n2430), .B(n15270), .ZN(n2427)
         );
  OAI22_X1 U1902 ( .A1(n14797), .A2(n15499), .B1(n3842), .B2(n14730), .ZN(
        n2430) );
  OAI221_X1 U1903 ( .B1(n9781), .B2(n14755), .C1(n9470), .C2(n14761), .A(n2443), .ZN(n2436) );
  AOI222_X1 U1904 ( .A1(n14837), .A2(n16089), .B1(n14824), .B2(n15543), .C1(
        n14782), .C2(n15580), .ZN(n2443) );
  OAI221_X1 U1905 ( .B1(n9401), .B2(n14762), .C1(n3697), .C2(n1471), .A(n2337), 
        .ZN(n2330) );
  AOI222_X1 U1906 ( .A1(n14747), .A2(n15851), .B1(n14726), .B2(n15865), .C1(
        n14825), .C2(n15746), .ZN(n2337) );
  INV_X1 U1907 ( .A(n2496), .ZN(n15295) );
  OAI221_X1 U1908 ( .B1(n14829), .B2(n3926), .C1(n1670), .C2(n3634), .A(n2497), 
        .ZN(n2496) );
  AOI221_X1 U1909 ( .B1(n15737), .B2(n14771), .C1(n14824), .C2(n9570), .A(
        Read_one_address[1]), .ZN(n2497) );
  INV_X1 U1910 ( .A(n2461), .ZN(n15296) );
  OAI221_X1 U1911 ( .B1(n14829), .B2(n3927), .C1(n1670), .C2(n3638), .A(n2462), 
        .ZN(n2461) );
  AOI221_X1 U1912 ( .B1(n15736), .B2(n14772), .C1(n14823), .C2(n9572), .A(
        Read_one_address[1]), .ZN(n2462) );
  OAI221_X1 U1913 ( .B1(n3287), .B2(n14813), .C1(n9363), .C2(n14718), .A(n2283), .ZN(n2275) );
  AOI21_X1 U1914 ( .B1(n14781), .B2(n15434), .A(n2154), .ZN(n2283) );
  OAI221_X1 U1915 ( .B1(n9862), .B2(n14762), .C1(n14829), .C2(n15374), .A(
        n2440), .ZN(n2439) );
  AOI22_X1 U1916 ( .A1(n14808), .A2(n16169), .B1(n14781), .B2(n15863), .ZN(
        n2440) );
  OAI221_X1 U1917 ( .B1(n3313), .B2(n14814), .C1(n9362), .C2(n14717), .A(n2153), .ZN(n2131) );
  AOI21_X1 U1918 ( .B1(n14782), .B2(n15433), .A(n2154), .ZN(n2153) );
  AOI211_X1 U1919 ( .C1(n14806), .C2(n16103), .A(n2498), .B(n2499), .ZN(n2495)
         );
  OAI21_X1 U1920 ( .B1(n3221), .B2(n14786), .A(n15277), .ZN(n2498) );
  AOI221_X1 U1921 ( .B1(n15291), .B2(n15423), .C1(n15292), .C2(n9607), .A(
        n1860), .ZN(n2499) );
  AOI211_X1 U1922 ( .C1(n14806), .C2(n16102), .A(n2463), .B(n2464), .ZN(n2460)
         );
  OAI21_X1 U1923 ( .B1(n3222), .B2(n14787), .A(n15277), .ZN(n2463) );
  AOI221_X1 U1924 ( .B1(n15291), .B2(n15421), .C1(n15292), .C2(n9609), .A(
        n1860), .ZN(n2464) );
  OAI221_X1 U1925 ( .B1(n1634), .B2(n15449), .C1(n3272), .C2(n14829), .A(n1657), .ZN(n2445) );
  OAI221_X1 U1926 ( .B1(n15912), .B2(n14797), .C1(n15921), .C2(n14761), .A(
        n2549), .ZN(n2547) );
  AOI22_X1 U1927 ( .A1(n14724), .A2(n3078), .B1(n14825), .B2(n3916), .ZN(n2549) );
  OAI221_X1 U1928 ( .B1(n2417), .B2(n2418), .C1(n2419), .C2(n2420), .A(n2322), 
        .ZN(n2416) );
  OAI221_X1 U1929 ( .B1(n9483), .B2(n14754), .C1(n3301), .C2(n14762), .A(n2422), .ZN(n2419) );
  OAI211_X1 U1930 ( .C1(n3194), .C2(n14828), .A(n15272), .B(n2421), .ZN(n2420)
         );
  OAI221_X1 U1931 ( .B1(n1634), .B2(n15448), .C1(n3273), .C2(n1471), .A(n1657), 
        .ZN(n2418) );
  AOI221_X1 U1932 ( .B1(n15285), .B2(n3868), .C1(n14848), .C2(Data_in[9]), .A(
        n2400), .ZN(n2399) );
  OAI222_X1 U1933 ( .A1(n16069), .A2(n1835), .B1(n15900), .B2(n1836), .C1(
        n3374), .C2(n1839), .ZN(n2400) );
  OAI221_X1 U1934 ( .B1(n16024), .B2(n2120), .C1(n14691), .C2(n14844), .A(
        n2122), .ZN(N983) );
  AOI222_X1 U1935 ( .A1(n1826), .A2(n9348), .B1(n2123), .B2(n14844), .C1(n1771), .C2(n3109), .ZN(n2122) );
  OAI221_X1 U1936 ( .B1(n2127), .B2(n2128), .C1(n2130), .C2(n2131), .A(n2137), 
        .ZN(n2123) );
  OAI221_X1 U1937 ( .B1(n9857), .B2(n14762), .C1(n9871), .C2(n1471), .A(n2157), 
        .ZN(n2127) );
  OAI221_X1 U1938 ( .B1(n3280), .B2(n14798), .C1(n3093), .C2(n14717), .A(n2338), .ZN(n2329) );
  AOI21_X1 U1939 ( .B1(n14781), .B2(n15694), .A(n1853), .ZN(n2338) );
  OAI221_X1 U1940 ( .B1(n9402), .B2(n14762), .C1(n3699), .C2(n14828), .A(n2284), .ZN(n2274) );
  AOI222_X1 U1941 ( .A1(n14807), .A2(n16248), .B1(n14748), .B2(n15910), .C1(
        n14742), .C2(n15752), .ZN(n2284) );
  OAI221_X1 U1942 ( .B1(n9398), .B2(n14762), .C1(n3698), .C2(n1471), .A(n2155), 
        .ZN(n2130) );
  AOI222_X1 U1943 ( .A1(n14807), .A2(n16247), .B1(n14748), .B2(n15908), .C1(
        n14742), .C2(n15751), .ZN(n2155) );
  OAI221_X1 U1944 ( .B1(n14749), .B2(n15478), .C1(n3944), .C2(n14730), .A(
        n2441), .ZN(n2438) );
  AOI221_X1 U1945 ( .B1(n14817), .B2(n15731), .C1(n14725), .C2(n16244), .A(
        n15271), .ZN(n2441) );
  OAI221_X1 U1946 ( .B1(n9656), .B2(n1652), .C1(n14797), .C2(n15349), .A(n1657), .ZN(n1715) );
  OAI221_X1 U1947 ( .B1(n9655), .B2(n1652), .C1(n14799), .C2(n15348), .A(n1657), .ZN(n1453) );
  OAI221_X1 U1948 ( .B1(n3305), .B2(n14828), .C1(n3850), .C2(n14730), .A(n1784), .ZN(n1776) );
  AOI21_X1 U1949 ( .B1(n14782), .B2(n15677), .A(n15270), .ZN(n1784) );
  OAI221_X1 U1950 ( .B1(n3867), .B2(n14718), .C1(n3659), .C2(n14812), .A(n1722), .ZN(n1703) );
  AOI21_X1 U1951 ( .B1(n14809), .B2(n16235), .A(n15270), .ZN(n1722) );
  OAI221_X1 U1952 ( .B1(n3644), .B2(n1670), .C1(n3660), .C2(n14812), .A(n1671), 
        .ZN(n1440) );
  AOI21_X1 U1953 ( .B1(n14809), .B2(n16234), .A(n15270), .ZN(n1671) );
  OAI221_X1 U1954 ( .B1(n3083), .B2(n14814), .C1(n9395), .C2(n14796), .A(n2264), .ZN(n2261) );
  AOI222_X1 U1955 ( .A1(n14783), .A2(n15509), .B1(n14726), .B2(n15842), .C1(
        n14742), .C2(n15607), .ZN(n2264) );
  OAI221_X1 U1956 ( .B1(n9528), .B2(n14718), .C1(n3088), .C2(n14813), .A(
        n15269), .ZN(n2259) );
  OAI221_X1 U1957 ( .B1(n9381), .B2(n14716), .C1(n3967), .C2(n14812), .A(
        n15269), .ZN(n1781) );
  OAI221_X1 U1958 ( .B1(n14749), .B2(n15398), .C1(n9411), .C2(n14761), .A(
        n2265), .ZN(n2258) );
  AOI22_X1 U1959 ( .A1(n14808), .A2(n16168), .B1(n14741), .B2(n16167), .ZN(
        n2265) );
  OAI221_X1 U1960 ( .B1(n9547), .B2(n14763), .C1(n9825), .C2(n1471), .A(n1783), 
        .ZN(n1780) );
  AOI22_X1 U1961 ( .A1(n14748), .A2(n15864), .B1(n14741), .B2(n16174), .ZN(
        n1783) );
  OAI22_X1 U1962 ( .A1(n3789), .A2(n14829), .B1(n14797), .B2(n15479), .ZN(
        n2210) );
  AOI221_X1 U1963 ( .B1(n14722), .B2(n9527), .C1(n14822), .C2(n15466), .A(
        n2350), .ZN(n2349) );
  OAI22_X1 U1964 ( .A1(n9582), .A2(n14751), .B1(n15992), .B2(n14795), .ZN(
        n2350) );
  OAI22_X1 U1965 ( .A1(n15784), .A2(n14730), .B1(n9442), .B2(n14759), .ZN(
        n2358) );
  OAI22_X1 U1966 ( .A1(n15785), .A2(n14730), .B1(n9440), .B2(n14759), .ZN(
        n2377) );
  OAI22_X1 U1967 ( .A1(n15783), .A2(n14729), .B1(n9891), .B2(n14760), .ZN(
        n2215) );
  OAI22_X1 U1968 ( .A1(n15782), .A2(n14729), .B1(n9441), .B2(n14759), .ZN(
        n2196) );
  AOI221_X1 U1969 ( .B1(n14782), .B2(n15389), .C1(n14839), .C2(n9868), .A(
        n2351), .ZN(n2348) );
  OAI22_X1 U1970 ( .A1(n16217), .A2(n14730), .B1(n3352), .B2(n14759), .ZN(
        n2351) );
  AOI221_X1 U1971 ( .B1(n14782), .B2(n15390), .C1(n14839), .C2(n9867), .A(
        n2370), .ZN(n2367) );
  OAI22_X1 U1972 ( .A1(n16218), .A2(n14730), .B1(n3351), .B2(n14759), .ZN(
        n2370) );
  OAI22_X1 U1973 ( .A1(n3255), .A2(n14785), .B1(n3298), .B2(n14760), .ZN(n2352) );
  OAI22_X1 U1974 ( .A1(n9820), .A2(n14829), .B1(n9883), .B2(n14759), .ZN(n2432) );
  OAI22_X1 U1975 ( .A1(n3254), .A2(n14784), .B1(n3286), .B2(n14759), .ZN(n2371) );
  OAI22_X1 U1976 ( .A1(n3257), .A2(n14784), .B1(n3875), .B2(n14759), .ZN(n2190) );
  OAI22_X1 U1977 ( .A1(n9473), .A2(n14760), .B1(n9498), .B2(n14752), .ZN(n1786) );
  OAI22_X1 U1978 ( .A1(n3903), .A2(n14784), .B1(n3246), .B2(n14795), .ZN(n1782) );
  OAI22_X1 U1979 ( .A1(n2544), .A2(n2545), .B1(n15278), .B2(n2546), .ZN(n2543)
         );
  OAI221_X1 U1980 ( .B1(n3345), .B2(n14718), .C1(n3853), .C2(n14812), .A(n2550), .ZN(n2545) );
  OAI221_X1 U1981 ( .B1(n3320), .B2(n14731), .C1(n9647), .C2(n14788), .A(n2551), .ZN(n2544) );
  AOI211_X1 U1982 ( .C1(n14836), .C2(n3202), .A(n2547), .B(n2548), .ZN(n2546)
         );
  OAI22_X1 U1983 ( .A1(n14762), .A2(n15354), .B1(n3805), .B2(n14751), .ZN(
        n1779) );
  AOI22_X1 U1984 ( .A1(n14738), .A2(n9640), .B1(n14783), .B2(n3886), .ZN(n2280) );
  AOI22_X1 U1985 ( .A1(n14739), .A2(n9641), .B1(n14783), .B2(n3914), .ZN(n2150) );
  OAI221_X1 U1986 ( .B1(n16026), .B2(n2120), .C1(n14670), .C2(n14844), .A(
        n2270), .ZN(N976) );
  AOI222_X1 U1987 ( .A1(n1826), .A2(n9350), .B1(n2271), .B2(n14844), .C1(n1771), .C2(n3108), .ZN(n2270) );
  OAI221_X1 U1988 ( .B1(n2272), .B2(n2273), .C1(n2274), .C2(n2275), .A(n2276), 
        .ZN(n2271) );
  OAI221_X1 U1989 ( .B1(n9856), .B2(n14763), .C1(n9870), .C2(n1471), .A(n2286), 
        .ZN(n2272) );
  OAI221_X1 U1990 ( .B1(n3288), .B2(n14798), .C1(n3933), .C2(n14787), .A(n2285), .ZN(n2273) );
  AOI21_X1 U1991 ( .B1(n3725), .B2(n14747), .A(n1853), .ZN(n2285) );
  OAI221_X1 U1992 ( .B1(n3315), .B2(n14798), .C1(n3833), .C2(n14787), .A(n2156), .ZN(n2128) );
  AOI21_X1 U1993 ( .B1(n3724), .B2(n14746), .A(n1853), .ZN(n2156) );
  INV_X1 U1994 ( .A(Read_one_address[4]), .ZN(n15347) );
  OAI211_X1 U1995 ( .C1(n3193), .C2(n14828), .A(n15272), .B(n2448), .ZN(n2447)
         );
  AOI22_X1 U1996 ( .A1(n14739), .A2(n16153), .B1(n14783), .B2(n16267), .ZN(
        n2448) );
  INV_X1 U1997 ( .A(Read_one_address[2]), .ZN(n15301) );
  OAI211_X1 U1998 ( .C1(n3817), .C2(n14797), .A(n15271), .B(n2442), .ZN(n2437)
         );
  AOI22_X1 U1999 ( .A1(n14738), .A2(n15647), .B1(n3640), .B2(n14719), .ZN(
        n2442) );
  OAI211_X1 U2000 ( .C1(n9378), .C2(n14797), .A(n15289), .B(n2336), .ZN(n2331)
         );
  AOI22_X1 U2001 ( .A1(n14738), .A2(n15541), .B1(n14781), .B2(n15432), .ZN(
        n2336) );
  OAI21_X1 U2002 ( .B1(n2509), .B2(n2510), .A(n2322), .ZN(n2508) );
  OAI221_X1 U2003 ( .B1(n9828), .B2(n14813), .C1(n9481), .C2(n14753), .A(n2511), .ZN(n2510) );
  OAI221_X1 U2004 ( .B1(n9644), .B2(n14789), .C1(n3378), .C2(n1471), .A(n2512), 
        .ZN(n2509) );
  AOI21_X1 U2005 ( .B1(n14740), .B2(n16087), .A(n15269), .ZN(n2511) );
  AOI221_X1 U2006 ( .B1(n3680), .B2(n15299), .C1(n14839), .C2(n16121), .A(
        n2224), .ZN(n2219) );
  OAI21_X1 U2007 ( .B1(n3104), .B2(n1652), .A(n2225), .ZN(n2224) );
  OAI221_X1 U2008 ( .B1(n14766), .B2(n16079), .C1(n15302), .C2(n16019), .A(
        n1650), .ZN(n2225) );
  AOI221_X1 U2009 ( .B1(n15299), .B2(n15685), .C1(n14838), .C2(n16123), .A(
        n2513), .ZN(n2507) );
  OAI21_X1 U2010 ( .B1(n3103), .B2(n1652), .A(n2514), .ZN(n2513) );
  OAI221_X1 U2011 ( .B1(n14766), .B2(n16082), .C1(n15302), .C2(n16022), .A(
        n1650), .ZN(n2514) );
  AOI221_X1 U2012 ( .B1(n3682), .B2(n15299), .C1(n14838), .C2(n16122), .A(
        n2295), .ZN(n2290) );
  OAI21_X1 U2013 ( .B1(n3105), .B2(n1652), .A(n2296), .ZN(n2295) );
  OAI221_X1 U2014 ( .B1(n14767), .B2(n16080), .C1(n15302), .C2(n16020), .A(
        n1650), .ZN(n2296) );
  AOI221_X1 U2015 ( .B1(n3681), .B2(n15299), .C1(n14841), .C2(n16120), .A(
        n2083), .ZN(n2071) );
  OAI21_X1 U2016 ( .B1(n3107), .B2(n1652), .A(n2084), .ZN(n2083) );
  OAI221_X1 U2017 ( .B1(n14766), .B2(n16078), .C1(n15302), .C2(n16018), .A(
        n1650), .ZN(n2084) );
  OAI211_X1 U2018 ( .C1(n3297), .C2(n1471), .A(n2180), .B(n2318), .ZN(n2315)
         );
  AOI22_X1 U2019 ( .A1(n14739), .A2(n15575), .B1(n14783), .B2(n15504), .ZN(
        n2318) );
  OAI211_X1 U2020 ( .C1(n3693), .C2(n1471), .A(n15289), .B(n2247), .ZN(n2244)
         );
  AOI22_X1 U2021 ( .A1(n14747), .A2(n15889), .B1(n14781), .B2(n15681), .ZN(
        n2247) );
  OAI211_X1 U2022 ( .C1(n3303), .C2(n1471), .A(n15289), .B(n2110), .ZN(n2107)
         );
  AOI22_X1 U2023 ( .A1(n14747), .A2(n15887), .B1(n14782), .B2(n15679), .ZN(
        n2110) );
  OAI211_X1 U2024 ( .C1(n3692), .C2(n1471), .A(n15289), .B(n2171), .ZN(n2168)
         );
  AOI22_X1 U2025 ( .A1(n14747), .A2(n15888), .B1(n14781), .B2(n15680), .ZN(
        n2171) );
  OAI211_X1 U2026 ( .C1(n3304), .C2(n1471), .A(n15289), .B(n1851), .ZN(n1848)
         );
  AOI22_X1 U2027 ( .A1(n14748), .A2(n15886), .B1(n14781), .B2(n15678), .ZN(
        n1851) );
  OAI211_X1 U2028 ( .C1(n3344), .C2(n1471), .A(n15289), .B(n2482), .ZN(n2479)
         );
  AOI22_X1 U2029 ( .A1(n14747), .A2(n15890), .B1(n14781), .B2(n15682), .ZN(
        n2482) );
  OAI211_X1 U2030 ( .C1(n3341), .C2(n1471), .A(n15289), .B(n2574), .ZN(n2571)
         );
  AOI22_X1 U2031 ( .A1(n14747), .A2(n15891), .B1(n14781), .B2(n15684), .ZN(
        n2574) );
  OAI21_X1 U2032 ( .B1(n3689), .B2(n14829), .A(n15276), .ZN(n2520) );
  OAI21_X1 U2033 ( .B1(n3688), .B2(n14829), .A(n15277), .ZN(n2557) );
  OAI21_X1 U2034 ( .B1(n3290), .B2(n14829), .A(n15274), .ZN(n2231) );
  OAI21_X1 U2035 ( .B1(n3808), .B2(n14828), .A(n15277), .ZN(n2538) );
  OAI21_X1 U2036 ( .B1(n3637), .B2(n14829), .A(n15276), .ZN(n2393) );
  OAI21_X1 U2037 ( .B1(n3289), .B2(n14829), .A(n15275), .ZN(n2302) );
  OAI21_X1 U2038 ( .B1(n3291), .B2(n14828), .A(n15274), .ZN(n2090) );
  OAI21_X1 U2039 ( .B1(n3292), .B2(n14828), .A(n15273), .ZN(n2055) );
  OAI21_X1 U2040 ( .B1(n3639), .B2(n14829), .A(n15274), .ZN(n1888) );
  OAI22_X1 U2041 ( .A1(n14646), .A2(n14845), .B1(n2414), .B2(n2415), .ZN(N968)
         );
  AOI221_X1 U2042 ( .B1(n2425), .B2(n2426), .C1(n2427), .C2(n2428), .A(n14618), 
        .ZN(n2414) );
  NAND2_X1 U2043 ( .A1(n2416), .A2(n14844), .ZN(n2415) );
  AOI221_X1 U2044 ( .B1(n3365), .B2(n14748), .C1(n14740), .C2(n16178), .A(
        n2432), .ZN(n2425) );
  OAI211_X1 U2045 ( .C1(n3955), .C2(n14718), .A(n14845), .B(n14619), .ZN(n2313) );
  OAI21_X1 U2046 ( .B1(n3953), .B2(n14811), .A(n15290), .ZN(n2353) );
  OAI21_X1 U2047 ( .B1(n3952), .B2(n14811), .A(n15290), .ZN(n2372) );
  OAI21_X1 U2048 ( .B1(n3865), .B2(n14829), .A(n1789), .ZN(n1787) );
  OAI21_X1 U2049 ( .B1(n16303), .B2(n1790), .A(n1792), .ZN(n1789) );
  OAI211_X1 U2050 ( .C1(n3293), .C2(n14730), .A(n14786), .B(n14845), .ZN(n1792) );
  NAND4_X1 U2051 ( .A1(n2340), .A2(n2341), .A3(n2342), .A4(n2343), .ZN(N972)
         );
  AOI22_X1 U2052 ( .A1(n15285), .A2(n3824), .B1(n14850), .B2(Data_in[12]), 
        .ZN(n2340) );
  AOI222_X1 U2053 ( .A1(n1826), .A2(n15381), .B1(n1771), .B2(n3129), .C1(n1793), .C2(n3061), .ZN(n2342) );
  AOI222_X1 U2054 ( .A1(n15288), .A2(n9837), .B1(n15287), .B2(n3181), .C1(
        n15286), .C2(n3330), .ZN(n2341) );
  NAND4_X1 U2055 ( .A1(n2359), .A2(n2360), .A3(n2361), .A4(n2362), .ZN(N971)
         );
  AOI22_X1 U2056 ( .A1(n15285), .A2(n3822), .B1(n14850), .B2(Data_in[11]), 
        .ZN(n2359) );
  AOI222_X1 U2057 ( .A1(n1826), .A2(n15382), .B1(n1771), .B2(n3128), .C1(n1793), .C2(n3060), .ZN(n2361) );
  AOI222_X1 U2058 ( .A1(n15288), .A2(n9836), .B1(n15287), .B2(n3180), .C1(
        n15286), .C2(n3328), .ZN(n2360) );
  NAND4_X1 U2059 ( .A1(n2197), .A2(n2198), .A3(n2199), .A4(n2200), .ZN(N980)
         );
  AOI22_X1 U2060 ( .A1(n15285), .A2(n9632), .B1(n14849), .B2(Data_in[20]), 
        .ZN(n2197) );
  AOI222_X1 U2061 ( .A1(n1826), .A2(n9790), .B1(n1771), .B2(n3106), .C1(n1793), 
        .C2(n9466), .ZN(n2199) );
  AOI222_X1 U2062 ( .A1(n15288), .A2(n15447), .B1(n15287), .B2(n3160), .C1(
        n15286), .C2(n9643), .ZN(n2198) );
  NAND4_X1 U2063 ( .A1(n2176), .A2(n2177), .A3(n2178), .A4(n2179), .ZN(N981)
         );
  AOI22_X1 U2064 ( .A1(n15285), .A2(n3135), .B1(n14849), .B2(Data_in[21]), 
        .ZN(n2176) );
  AOI222_X1 U2065 ( .A1(n1826), .A2(n15380), .B1(n1771), .B2(n3130), .C1(n1793), .C2(n3062), .ZN(n2178) );
  AOI222_X1 U2066 ( .A1(n15288), .A2(n9835), .B1(n15287), .B2(n3182), .C1(
        n15286), .C2(n3332), .ZN(n2177) );
  NAND4_X1 U2067 ( .A1(n1767), .A2(n1768), .A3(n1769), .A4(n1770), .ZN(N989)
         );
  AOI22_X1 U2068 ( .A1(n1793), .A2(n3339), .B1(n1826), .B2(n9347), .ZN(n1769)
         );
  AOI22_X1 U2069 ( .A1(n15285), .A2(n3178), .B1(n14849), .B2(Data_in[29]), 
        .ZN(n1767) );
  AOI222_X1 U2070 ( .A1(n15288), .A2(n15446), .B1(n15287), .B2(n3641), .C1(
        n15286), .C2(n3299), .ZN(n1768) );
  INV_X1 U2071 ( .A(Read_one_address[3]), .ZN(n15303) );
  NAND4_X1 U2072 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(N969)
         );
  NAND4_X1 U2073 ( .A1(n15278), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2397)
         );
  AOI222_X1 U2074 ( .A1(n1826), .A2(n9492), .B1(n1771), .B2(n3059), .C1(n1793), 
        .C2(n3948), .ZN(n2398) );
  AOI22_X1 U2075 ( .A1(n2406), .A2(n2407), .B1(n2408), .B2(n2409), .ZN(n2396)
         );
  AOI222_X1 U2076 ( .A1(n1826), .A2(n9495), .B1(n1771), .B2(n3069), .C1(n1793), 
        .C2(n3957), .ZN(n2305) );
  AOI21_X1 U2077 ( .B1(n2309), .B2(n2310), .A(n2311), .ZN(n2306) );
  AOI221_X1 U2078 ( .B1(n15285), .B2(n9627), .C1(n14849), .C2(Data_in[14]), 
        .A(n2308), .ZN(n2307) );
  AOI222_X1 U2079 ( .A1(n1826), .A2(n9493), .B1(n1771), .B2(n3057), .C1(n1793), 
        .C2(n3212), .ZN(n2487) );
  AOI221_X1 U2080 ( .B1(n15285), .B2(n9629), .C1(n14847), .C2(Data_in[4]), .A(
        n2490), .ZN(n2489) );
  AOI222_X1 U2081 ( .A1(n2491), .A2(n2492), .B1(n2493), .B2(n2494), .C1(n2495), 
        .C2(n15295), .ZN(n2488) );
  AOI222_X1 U2082 ( .A1(n1826), .A2(n9494), .B1(n1771), .B2(n3058), .C1(n1793), 
        .C2(n3231), .ZN(n2452) );
  AOI221_X1 U2083 ( .B1(n15285), .B2(n9630), .C1(n14847), .C2(Data_in[6]), .A(
        n2455), .ZN(n2454) );
  AOI222_X1 U2084 ( .A1(n2456), .A2(n2457), .B1(n2458), .B2(n2459), .C1(n2460), 
        .C2(n15296), .ZN(n2453) );
  BUF_X1 U2085 ( .A(n1670), .Z(n14716) );
  NAND2_X1 U2086 ( .A1(n15300), .A2(Read_one_address[4]), .ZN(n1670) );
  BUF_X1 U2087 ( .A(n1662), .Z(n14758) );
  BUF_X1 U2088 ( .A(n1656), .Z(n14794) );
  NAND2_X1 U2089 ( .A1(n2355), .A2(n2356), .ZN(n2344) );
  AOI221_X1 U2090 ( .B1(n14721), .B2(n15377), .C1(n14822), .C2(n3959), .A(
        n2357), .ZN(n2356) );
  AOI221_X1 U2091 ( .B1(n14782), .B2(n3977), .C1(n14838), .C2(n3110), .A(n2358), .ZN(n2355) );
  OAI22_X1 U2092 ( .A1(n3347), .A2(n14751), .B1(n16312), .B2(n14796), .ZN(
        n2357) );
  NAND2_X1 U2093 ( .A1(n2374), .A2(n2375), .ZN(n2363) );
  AOI221_X1 U2094 ( .B1(n14721), .B2(n15378), .C1(n14823), .C2(n3958), .A(
        n2376), .ZN(n2375) );
  AOI221_X1 U2095 ( .B1(n14781), .B2(n3976), .C1(n14840), .C2(n3114), .A(n2377), .ZN(n2374) );
  OAI22_X1 U2096 ( .A1(n3346), .A2(n14751), .B1(n16313), .B2(n14795), .ZN(
        n2376) );
  NAND2_X1 U2097 ( .A1(n2212), .A2(n2213), .ZN(n2201) );
  AOI221_X1 U2098 ( .B1(n14720), .B2(n9524), .C1(n14820), .C2(n3089), .A(n2214), .ZN(n2213) );
  AOI221_X1 U2099 ( .B1(n14782), .B2(n3053), .C1(n14839), .C2(n3123), .A(n2215), .ZN(n2212) );
  OAI22_X1 U2100 ( .A1(n15905), .A2(n14750), .B1(n16199), .B2(n14796), .ZN(
        n2214) );
  NAND2_X1 U2101 ( .A1(n2193), .A2(n2194), .ZN(n2181) );
  AOI221_X1 U2102 ( .B1(n14720), .B2(n15376), .C1(n14820), .C2(n3960), .A(
        n2195), .ZN(n2194) );
  AOI221_X1 U2103 ( .B1(n14782), .B2(n3978), .C1(n14840), .C2(n3115), .A(n2196), .ZN(n2193) );
  OAI22_X1 U2104 ( .A1(n3348), .A2(n14749), .B1(n16311), .B2(n14796), .ZN(
        n2195) );
  AOI22_X1 U2105 ( .A1(n1793), .A2(n3082), .B1(n1826), .B2(n9793), .ZN(n2234)
         );
  AOI221_X1 U2106 ( .B1(n15285), .B2(n3112), .C1(n14848), .C2(Data_in[18]), 
        .A(n2237), .ZN(n2236) );
  AOI222_X1 U2107 ( .A1(n1771), .A2(n3074), .B1(n2238), .B2(n2239), .C1(n2240), 
        .C2(n14845), .ZN(n2235) );
  AOI22_X1 U2108 ( .A1(n1793), .A2(n3087), .B1(n1826), .B2(n9795), .ZN(n2095)
         );
  AOI221_X1 U2109 ( .B1(n15285), .B2(n3116), .C1(n14846), .C2(Data_in[24]), 
        .A(n2098), .ZN(n2097) );
  AOI222_X1 U2110 ( .A1(n1771), .A2(n3076), .B1(n2099), .B2(n2100), .C1(n2101), 
        .C2(n14845), .ZN(n2096) );
  AOI22_X1 U2111 ( .A1(n1793), .A2(n3086), .B1(n1826), .B2(n9794), .ZN(n2158)
         );
  AOI221_X1 U2112 ( .B1(n15285), .B2(n3113), .C1(n14847), .C2(Data_in[22]), 
        .A(n2161), .ZN(n2160) );
  AOI222_X1 U2113 ( .A1(n1771), .A2(n3075), .B1(n2162), .B2(n2163), .C1(n2164), 
        .C2(n14845), .ZN(n2159) );
  AOI22_X1 U2114 ( .A1(n1793), .A2(n3081), .B1(n1826), .B2(n9792), .ZN(n2469)
         );
  AOI221_X1 U2115 ( .B1(n15285), .B2(n3111), .C1(n14847), .C2(Data_in[5]), .A(
        n2472), .ZN(n2471) );
  AOI222_X1 U2116 ( .A1(n1771), .A2(n3072), .B1(n2473), .B2(n2474), .C1(n2475), 
        .C2(n14845), .ZN(n2470) );
  AOI22_X1 U2117 ( .A1(n1793), .A2(n3080), .B1(n1826), .B2(n9791), .ZN(n2560)
         );
  AOI221_X1 U2118 ( .B1(n15285), .B2(n3098), .C1(n14846), .C2(Data_in[0]), .A(
        n2563), .ZN(n2562) );
  AOI222_X1 U2119 ( .A1(n1771), .A2(n3071), .B1(n2565), .B2(n2566), .C1(n2567), 
        .C2(n14844), .ZN(n2561) );
  AOI22_X1 U2120 ( .A1(n1793), .A2(n3092), .B1(n1826), .B2(n9796), .ZN(n1828)
         );
  AOI221_X1 U2121 ( .B1(n15285), .B2(n3127), .C1(n14846), .C2(Data_in[28]), 
        .A(n1832), .ZN(n1831) );
  AOI222_X1 U2122 ( .A1(n1771), .A2(n3077), .B1(n1840), .B2(n1841), .C1(n1842), 
        .C2(n14845), .ZN(n1830) );
  NAND2_X1 U2123 ( .A1(n15299), .A2(Read_one_address[3]), .ZN(n1658) );
  AOI22_X1 U2124 ( .A1(n1793), .A2(n3302), .B1(n1826), .B2(n9789), .ZN(n2252)
         );
  AOI221_X1 U2125 ( .B1(n15285), .B2(n3140), .C1(n14848), .C2(Data_in[17]), 
        .A(n2255), .ZN(n2254) );
  AOI222_X1 U2126 ( .A1(n1771), .A2(n3073), .B1(n2256), .B2(n15297), .C1(
        n15293), .C2(n2257), .ZN(n2253) );
  AOI22_X1 U2127 ( .A1(n1826), .A2(n9349), .B1(n15287), .B2(n3700), .ZN(n2323)
         );
  AOI221_X1 U2128 ( .B1(n15285), .B2(n3279), .C1(n14848), .C2(Data_in[13]), 
        .A(n2326), .ZN(n2325) );
  AOI222_X1 U2129 ( .A1(n1793), .A2(n9462), .B1(n2327), .B2(n14844), .C1(n1771), .C2(n3099), .ZN(n2324) );
  BUF_X1 U2130 ( .A(n1471), .Z(n14828) );
  INV_X1 U2131 ( .A(n2266), .ZN(n15297) );
  OAI221_X1 U2132 ( .B1(n14829), .B2(n3928), .C1(n1670), .C2(n3851), .A(n2267), 
        .ZN(n2266) );
  AOI221_X1 U2133 ( .B1(n15735), .B2(n14772), .C1(n14821), .C2(n9571), .A(
        Read_one_address[1]), .ZN(n2267) );
  OAI21_X1 U2134 ( .B1(n14643), .B2(n14845), .A(n2433), .ZN(N967) );
  OAI221_X1 U2135 ( .B1(n2436), .B2(n2437), .C1(n2438), .C2(n2439), .A(
        Read_one_address[1]), .ZN(n2435) );
  OAI221_X1 U2136 ( .B1(n2444), .B2(n2445), .C1(n2446), .C2(n2447), .A(n2322), 
        .ZN(n2434) );
  NAND2_X1 U2137 ( .A1(Read_one_address[1]), .A2(n14844), .ZN(n2322) );
  NAND2_X1 U2138 ( .A1(Read_one_address[1]), .A2(n15270), .ZN(n1853) );
  OAI222_X1 U2139 ( .A1(n9335), .A2(n14756), .B1(n3271), .B2(n14816), .C1(
        n9365), .C2(n14763), .ZN(n1690) );
  AOI221_X1 U2140 ( .B1(n14836), .B2(n16043), .C1(n14740), .C2(n15577), .A(
        n2465), .ZN(n2459) );
  OAI222_X1 U2141 ( .A1(n9479), .A2(n14799), .B1(n3864), .B2(n14816), .C1(
        n9399), .C2(n14763), .ZN(n2465) );
  AOI221_X1 U2142 ( .B1(n14767), .B2(n15715), .C1(n14838), .C2(n15795), .A(
        n2320), .ZN(n2310) );
  OAI221_X1 U2143 ( .B1(n3275), .B2(n14797), .C1(n14756), .C2(n15450), .A(
        n15269), .ZN(n2320) );
  AOI221_X1 U2144 ( .B1(n15299), .B2(n15444), .C1(n14840), .C2(n15930), .A(
        n2531), .ZN(n2526) );
  OAI22_X1 U2145 ( .A1(n14797), .A2(n15353), .B1(n9612), .B2(n1652), .ZN(n2531) );
  AOI221_X1 U2146 ( .B1(n15299), .B2(n15443), .C1(n14837), .C2(n15929), .A(
        n2386), .ZN(n2381) );
  OAI22_X1 U2147 ( .A1(n14797), .A2(n15352), .B1(n9613), .B2(n1652), .ZN(n2386) );
  AOI221_X1 U2148 ( .B1(n14767), .B2(n15563), .C1(n14739), .C2(n16104), .A(
        n2404), .ZN(n2403) );
  OAI221_X1 U2149 ( .B1(n9872), .B2(n14813), .C1(n14799), .C2(n15481), .A(
        n14618), .ZN(n2404) );
  OAI221_X1 U2150 ( .B1(n9482), .B2(n14755), .C1(n3300), .C2(n14761), .A(n2449), .ZN(n2446) );
  AOI222_X1 U2151 ( .A1(n14807), .A2(n16150), .B1(n14726), .B2(n15954), .C1(
        n14825), .C2(n15670), .ZN(n2449) );
  NAND2_X1 U2152 ( .A1(Read_one_address[1]), .A2(n15271), .ZN(n2154) );
  NOR2_X1 U2153 ( .A1(n15272), .A2(Read_one_address[1]), .ZN(n2148) );
  AOI21_X1 U2154 ( .B1(n3657), .B2(n14765), .A(n1853), .ZN(n2248) );
  AOI21_X1 U2155 ( .B1(n3656), .B2(n14764), .A(n1853), .ZN(n2111) );
  AOI21_X1 U2156 ( .B1(n3653), .B2(n14764), .A(n1853), .ZN(n2172) );
  AOI21_X1 U2157 ( .B1(n3658), .B2(n14765), .A(n1853), .ZN(n2483) );
  AOI21_X1 U2158 ( .B1(n3655), .B2(n14765), .A(n1853), .ZN(n2575) );
  AOI21_X1 U2159 ( .B1(n3654), .B2(n14764), .A(n1853), .ZN(n1852) );
  INV_X1 U2160 ( .A(Read_one_address[1]), .ZN(n15294) );
  OAI211_X1 U2161 ( .C1(n9546), .C2(n14813), .A(n14845), .B(n14619), .ZN(n2209) );
  OAI21_X1 U2162 ( .B1(n3147), .B2(n14846), .A(n2405), .ZN(n2401) );
  OAI21_X1 U2163 ( .B1(n3892), .B2(n14811), .A(n15290), .ZN(n2191) );
  BUF_X1 U2164 ( .A(Read_one_address[0]), .Z(n15267) );
  BUF_X1 U2165 ( .A(Read_one_address[0]), .Z(n15266) );
  BUF_X1 U2166 ( .A(Read_one_address[0]), .Z(n15268) );
  NOR3_X1 U2167 ( .A1(n15283), .A2(Read_two_address[4]), .A3(n15282), .ZN(
        n3029) );
  NOR3_X1 U2168 ( .A1(n15282), .A2(Read_two_address[3]), .A3(n15284), .ZN(
        n3033) );
  NOR3_X1 U2169 ( .A1(Read_two_address[2]), .A2(Read_two_address[4]), .A3(
        n15283), .ZN(n3026) );
  NOR3_X1 U2170 ( .A1(n15283), .A2(Read_two_address[2]), .A3(n15284), .ZN(
        n3028) );
  NOR3_X1 U2171 ( .A1(Read_two_address[2]), .A2(Read_two_address[3]), .A3(
        n15284), .ZN(n3034) );
  NOR3_X1 U2172 ( .A1(Read_two_address[3]), .A2(Read_two_address[4]), .A3(
        n15282), .ZN(n3027) );
  NOR3_X1 U2173 ( .A1(Read_two_address[3]), .A2(Read_two_address[4]), .A3(
        Read_two_address[2]), .ZN(n3031) );
  OAI221_X1 U2174 ( .B1(n9570), .B2(n14946), .C1(n15737), .C2(n14943), .A(
        n1274), .ZN(n1272) );
  AOI22_X1 U2175 ( .A1(n14940), .A2(n9607), .B1(n14935), .B2(n3221), .ZN(n1274) );
  OAI221_X1 U2176 ( .B1(n9572), .B2(n14946), .C1(n15736), .C2(n14943), .A(
        n1136), .ZN(n1133) );
  AOI22_X1 U2177 ( .A1(n14940), .A2(n9609), .B1(n14935), .B2(n3222), .ZN(n1136) );
  OAI221_X1 U2178 ( .B1(n9571), .B2(n14944), .C1(n15735), .C2(n14941), .A(
        n2844), .ZN(n2843) );
  AOI22_X1 U2179 ( .A1(n14938), .A2(n9608), .B1(n14936), .B2(n3223), .ZN(n2844) );
  OAI221_X1 U2180 ( .B1(n9733), .B2(n14898), .C1(n15444), .C2(n14895), .A(
        n1332), .ZN(n1329) );
  AOI22_X1 U2181 ( .A1(n14892), .A2(n3095), .B1(n14889), .B2(Data_in[2]), .ZN(
        n1332) );
  OAI221_X1 U2182 ( .B1(n9732), .B2(n14896), .C1(n15443), .C2(n14893), .A(
        n2978), .ZN(n2977) );
  AOI22_X1 U2183 ( .A1(n14890), .A2(n3843), .B1(n14887), .B2(Data_in[10]), 
        .ZN(n2978) );
  OAI221_X1 U2184 ( .B1(n9736), .B2(n14897), .C1(n15442), .C2(n14894), .A(
        n2690), .ZN(n2689) );
  AOI22_X1 U2185 ( .A1(n14891), .A2(n3848), .B1(n14888), .B2(Data_in[26]), 
        .ZN(n2690) );
  OAI221_X1 U2186 ( .B1(n9740), .B2(n14897), .C1(n15441), .C2(n14894), .A(
        n2672), .ZN(n2671) );
  AOI22_X1 U2187 ( .A1(n14891), .A2(n3849), .B1(n14889), .B2(Data_in[27]), 
        .ZN(n2672) );
  OAI221_X1 U2188 ( .B1(n9737), .B2(n14897), .C1(n15440), .C2(n14894), .A(
        n2618), .ZN(n2617) );
  AOI22_X1 U2189 ( .A1(n14891), .A2(n3939), .B1(n14889), .B2(Data_in[30]), 
        .ZN(n2618) );
  OAI221_X1 U2190 ( .B1(n9738), .B2(n14898), .C1(n15439), .C2(n14895), .A(
        n2600), .ZN(n2599) );
  AOI22_X1 U2191 ( .A1(n14892), .A2(n3832), .B1(n14889), .B2(Data_in[31]), 
        .ZN(n2600) );
  OAI221_X1 U2192 ( .B1(n9734), .B2(n14896), .C1(n3682), .C2(n14893), .A(n2888), .ZN(n2887) );
  AOI22_X1 U2193 ( .A1(n14890), .A2(n3844), .B1(n14888), .B2(Data_in[15]), 
        .ZN(n2888) );
  OAI221_X1 U2194 ( .B1(n9735), .B2(n14897), .C1(n3680), .C2(n14894), .A(n2816), .ZN(n2815) );
  AOI22_X1 U2195 ( .A1(n14891), .A2(n3845), .B1(n14888), .B2(Data_in[19]), 
        .ZN(n2816) );
  OAI221_X1 U2196 ( .B1(n9739), .B2(n14897), .C1(n3681), .C2(n14894), .A(n2708), .ZN(n2707) );
  AOI22_X1 U2197 ( .A1(n14891), .A2(n3847), .B1(n14888), .B2(Data_in[25]), 
        .ZN(n2708) );
  OAI221_X1 U2198 ( .B1(n15530), .B2(n14946), .C1(n15557), .C2(n14943), .A(
        n1420), .ZN(n1418) );
  AOI22_X1 U2199 ( .A1(n14940), .A2(n9602), .B1(n14935), .B2(n3712), .ZN(n1420) );
  OAI221_X1 U2200 ( .B1(n15904), .B2(n14898), .C1(n15614), .C2(n14895), .A(
        n1432), .ZN(n1429) );
  AOI22_X1 U2201 ( .A1(n14892), .A2(n3666), .B1(n14889), .B2(Data_in[0]), .ZN(
        n1432) );
  OAI221_X1 U2202 ( .B1(n15579), .B2(n14946), .C1(n15532), .C2(n14943), .A(
        n1345), .ZN(n1344) );
  AOI22_X1 U2203 ( .A1(n14940), .A2(n3320), .B1(n14935), .B2(n9647), .ZN(n1345) );
  OAI221_X1 U2204 ( .B1(n15912), .B2(n14898), .C1(n15613), .C2(n14895), .A(
        n1398), .ZN(n1397) );
  AOI22_X1 U2205 ( .A1(n14892), .A2(n3684), .B1(n14889), .B2(Data_in[1]), .ZN(
        n1398) );
  OAI221_X1 U2206 ( .B1(n15503), .B2(n14946), .C1(n15637), .C2(n14943), .A(
        n1314), .ZN(n1313) );
  AOI22_X1 U2207 ( .A1(n14940), .A2(n9659), .B1(n14935), .B2(n3213), .ZN(n1314) );
  OAI221_X1 U2208 ( .B1(n15583), .B2(n14946), .C1(n15508), .C2(n14943), .A(
        n1295), .ZN(n1292) );
  AOI22_X1 U2209 ( .A1(n14940), .A2(n3283), .B1(n14935), .B2(n9644), .ZN(n1295) );
  OAI221_X1 U2210 ( .B1(n15789), .B2(n14898), .C1(n15685), .C2(n14895), .A(
        n1304), .ZN(n1302) );
  AOI22_X1 U2211 ( .A1(n14892), .A2(n3840), .B1(n14889), .B2(Data_in[3]), .ZN(
        n1304) );
  OAI221_X1 U2212 ( .B1(n15903), .B2(n14898), .C1(n3372), .C2(n14895), .A(
        n1282), .ZN(n1281) );
  AOI22_X1 U2213 ( .A1(n14892), .A2(n3696), .B1(n14889), .B2(Data_in[4]), .ZN(
        n1282) );
  OAI221_X1 U2214 ( .B1(n15529), .B2(n14946), .C1(n15556), .C2(n14943), .A(
        n1227), .ZN(n1224) );
  AOI22_X1 U2215 ( .A1(n14940), .A2(n9601), .B1(n14935), .B2(n3232), .ZN(n1227) );
  OAI221_X1 U2216 ( .B1(n15902), .B2(n14898), .C1(n15612), .C2(n14895), .A(
        n1250), .ZN(n1241) );
  AOI22_X1 U2217 ( .A1(n14892), .A2(n3818), .B1(n14887), .B2(Data_in[5]), .ZN(
        n1250) );
  OAI221_X1 U2218 ( .B1(n15901), .B2(n14898), .C1(n3373), .C2(n14895), .A(
        n1162), .ZN(n1159) );
  AOI22_X1 U2219 ( .A1(n14892), .A2(n3831), .B1(n14888), .B2(Data_in[6]), .ZN(
        n1162) );
  OAI221_X1 U2220 ( .B1(n15520), .B2(n14946), .C1(n15430), .C2(n14943), .A(
        n2592), .ZN(n2591) );
  AOI22_X1 U2221 ( .A1(n14940), .A2(n3325), .B1(n14935), .B2(n3322), .ZN(n2592) );
  OAI221_X1 U2222 ( .B1(n15670), .B2(n14944), .C1(n15619), .C2(n14941), .A(
        n3024), .ZN(n3023) );
  AOI22_X1 U2223 ( .A1(n14938), .A2(n3284), .B1(n14937), .B2(n9645), .ZN(n3024) );
  OAI221_X1 U2224 ( .B1(n15788), .B2(n14896), .C1(n9502), .C2(n14893), .A(
        n3044), .ZN(n3043) );
  AOI22_X1 U2225 ( .A1(n14890), .A2(n3841), .B1(n14887), .B2(Data_in[7]), .ZN(
        n3044) );
  OAI221_X1 U2226 ( .B1(n15669), .B2(n14944), .C1(n15618), .C2(n14941), .A(
        n3006), .ZN(n3005) );
  AOI22_X1 U2227 ( .A1(n14938), .A2(n3285), .B1(n14937), .B2(n9646), .ZN(n3006) );
  OAI221_X1 U2228 ( .B1(n15787), .B2(n14896), .C1(n9503), .C2(n14893), .A(
        n3014), .ZN(n3013) );
  AOI22_X1 U2229 ( .A1(n14890), .A2(n3842), .B1(n14887), .B2(Data_in[8]), .ZN(
        n3014) );
  OAI221_X1 U2230 ( .B1(n15651), .B2(n14944), .C1(n15563), .C2(n14941), .A(
        n2988), .ZN(n2987) );
  AOI22_X1 U2231 ( .A1(n14938), .A2(n3673), .B1(n14937), .B2(n3260), .ZN(n2988) );
  OAI221_X1 U2232 ( .B1(n15900), .B2(n14896), .C1(n3374), .C2(n14893), .A(
        n2996), .ZN(n2995) );
  AOI22_X1 U2233 ( .A1(n14890), .A2(n3876), .B1(n14887), .B2(Data_in[9]), .ZN(
        n2996) );
  OAI221_X1 U2234 ( .B1(n15502), .B2(n14944), .C1(n15636), .C2(n14941), .A(
        n2970), .ZN(n2969) );
  AOI22_X1 U2235 ( .A1(n14938), .A2(n9660), .B1(n14937), .B2(n3214), .ZN(n2970) );
  OAI221_X1 U2236 ( .B1(n15513), .B2(n14944), .C1(n15745), .C2(n14941), .A(
        n2952), .ZN(n2951) );
  AOI22_X1 U2237 ( .A1(n14938), .A2(n9605), .B1(n14937), .B2(n3254), .ZN(n2952) );
  OAI221_X1 U2238 ( .B1(n15916), .B2(n14896), .C1(n15734), .C2(n14893), .A(
        n2960), .ZN(n2959) );
  AOI22_X1 U2239 ( .A1(n14890), .A2(n3895), .B1(n14887), .B2(Data_in[11]), 
        .ZN(n2960) );
  OAI221_X1 U2241 ( .B1(n15512), .B2(n14944), .C1(n15744), .C2(n14941), .A(
        n2934), .ZN(n2933) );
  AOI22_X1 U2242 ( .A1(n14938), .A2(n9604), .B1(n14937), .B2(n3255), .ZN(n2934) );
  OAI221_X1 U2243 ( .B1(n15915), .B2(n14896), .C1(n15733), .C2(n14893), .A(
        n2942), .ZN(n2941) );
  AOI22_X1 U2244 ( .A1(n14890), .A2(n3896), .B1(n14887), .B2(Data_in[12]), 
        .ZN(n2942) );
  OAI221_X1 U2245 ( .B1(n15581), .B2(n14944), .C1(n15587), .C2(n14941), .A(
        n2916), .ZN(n2915) );
  AOI22_X1 U2246 ( .A1(n14938), .A2(n3716), .B1(n14937), .B2(n3267), .ZN(n2916) );
  OAI221_X1 U2247 ( .B1(n15899), .B2(n14896), .C1(n15633), .C2(n14893), .A(
        n2924), .ZN(n2923) );
  AOI22_X1 U2248 ( .A1(n14890), .A2(n3877), .B1(n14887), .B2(Data_in[13]), 
        .ZN(n2924) );
  OAI221_X1 U2249 ( .B1(n15582), .B2(n14944), .C1(n9450), .C2(n14941), .A(
        n2898), .ZN(n2897) );
  AOI22_X1 U2250 ( .A1(n14938), .A2(n15482), .B1(n14937), .B2(n3256), .ZN(
        n2898) );
  OAI221_X1 U2251 ( .B1(n15898), .B2(n14896), .C1(n3375), .C2(n14893), .A(
        n2906), .ZN(n2905) );
  AOI22_X1 U2252 ( .A1(n14890), .A2(n3880), .B1(n14887), .B2(Data_in[14]), 
        .ZN(n2906) );
  OAI221_X1 U2253 ( .B1(n15528), .B2(n14944), .C1(n15617), .C2(n14941), .A(
        n2880), .ZN(n2879) );
  AOI22_X1 U2254 ( .A1(n14938), .A2(n3678), .B1(n14936), .B2(n3677), .ZN(n2880) );
  OAI221_X1 U2255 ( .B1(n15586), .B2(n14944), .C1(n15555), .C2(n14941), .A(
        n2862), .ZN(n2861) );
  AOI22_X1 U2256 ( .A1(n14938), .A2(n3720), .B1(n14936), .B2(n3665), .ZN(n2862) );
  OAI221_X1 U2257 ( .B1(n15918), .B2(n14896), .C1(n15496), .C2(n14893), .A(
        n2870), .ZN(n2869) );
  AOI22_X1 U2258 ( .A1(n14890), .A2(n3900), .B1(n14888), .B2(Data_in[16]), 
        .ZN(n2870) );
  OAI221_X1 U2259 ( .B1(n15897), .B2(n14896), .C1(n3379), .C2(n14893), .A(
        n2852), .ZN(n2851) );
  AOI22_X1 U2260 ( .A1(n14890), .A2(n3146), .B1(n14888), .B2(Data_in[17]), 
        .ZN(n2852) );
  OAI221_X1 U2261 ( .B1(n15527), .B2(n14944), .C1(n15554), .C2(n14941), .A(
        n2826), .ZN(n2825) );
  AOI22_X1 U2262 ( .A1(n14938), .A2(n9598), .B1(n14936), .B2(n3233), .ZN(n2826) );
  OAI221_X1 U2263 ( .B1(n15896), .B2(n14896), .C1(n15611), .C2(n14893), .A(
        n2834), .ZN(n2833) );
  AOI22_X1 U2264 ( .A1(n14890), .A2(n3889), .B1(n14888), .B2(Data_in[18]), 
        .ZN(n2834) );
  OAI221_X1 U2265 ( .B1(n15526), .B2(n14945), .C1(n15616), .C2(n14942), .A(
        n2808), .ZN(n2807) );
  AOI22_X1 U2266 ( .A1(n14939), .A2(n3312), .B1(n14936), .B2(n3261), .ZN(n2808) );
  OAI221_X1 U2267 ( .B1(n15585), .B2(n14945), .C1(n15456), .C2(n14942), .A(
        n2790), .ZN(n2789) );
  AOI22_X1 U2268 ( .A1(n14939), .A2(n3703), .B1(n14936), .B2(n3269), .ZN(n2790) );
  OAI221_X1 U2269 ( .B1(n15914), .B2(n14897), .C1(n3382), .C2(n14894), .A(
        n2798), .ZN(n2797) );
  AOI22_X1 U2270 ( .A1(n14891), .A2(n3846), .B1(n14888), .B2(Data_in[20]), 
        .ZN(n2798) );
  OAI221_X1 U2271 ( .B1(n15511), .B2(n14945), .C1(n15743), .C2(n14942), .A(
        n2772), .ZN(n2771) );
  AOI22_X1 U2272 ( .A1(n14939), .A2(n9606), .B1(n14936), .B2(n3257), .ZN(n2772) );
  OAI221_X1 U2273 ( .B1(n15913), .B2(n14897), .C1(n15732), .C2(n14894), .A(
        n2780), .ZN(n2779) );
  AOI22_X1 U2274 ( .A1(n14891), .A2(n3897), .B1(n14888), .B2(Data_in[21]), 
        .ZN(n2780) );
  OAI221_X1 U2275 ( .B1(n15525), .B2(n14945), .C1(n15553), .C2(n14942), .A(
        n2754), .ZN(n2753) );
  AOI22_X1 U2276 ( .A1(n14939), .A2(n9600), .B1(n14936), .B2(n3234), .ZN(n2754) );
  OAI221_X1 U2277 ( .B1(n15895), .B2(n14897), .C1(n15610), .C2(n14894), .A(
        n2762), .ZN(n2761) );
  AOI22_X1 U2278 ( .A1(n14891), .A2(n3899), .B1(n14888), .B2(Data_in[22]), 
        .ZN(n2762) );
  OAI221_X1 U2279 ( .B1(n15584), .B2(n14945), .C1(n15552), .C2(n14942), .A(
        n2736), .ZN(n2735) );
  AOI22_X1 U2280 ( .A1(n14939), .A2(n3718), .B1(n14936), .B2(n3652), .ZN(n2736) );
  OAI221_X1 U2281 ( .B1(n15917), .B2(n14897), .C1(n15495), .C2(n14894), .A(
        n2744), .ZN(n2743) );
  AOI22_X1 U2282 ( .A1(n14891), .A2(n3898), .B1(n14888), .B2(Data_in[23]), 
        .ZN(n2744) );
  OAI221_X1 U2283 ( .B1(n15524), .B2(n14945), .C1(n15551), .C2(n14942), .A(
        n2718), .ZN(n2717) );
  AOI22_X1 U2284 ( .A1(n14939), .A2(n9599), .B1(n14936), .B2(n3235), .ZN(n2718) );
  OAI221_X1 U2285 ( .B1(n15894), .B2(n14897), .C1(n15609), .C2(n14894), .A(
        n2726), .ZN(n2725) );
  AOI22_X1 U2286 ( .A1(n14891), .A2(n3919), .B1(n14888), .B2(Data_in[24]), 
        .ZN(n2726) );
  OAI221_X1 U2287 ( .B1(n15523), .B2(n14945), .C1(n15615), .C2(n14942), .A(
        n2700), .ZN(n2699) );
  AOI22_X1 U2288 ( .A1(n14939), .A2(n3676), .B1(n14936), .B2(n3675), .ZN(n2700) );
  OAI221_X1 U2289 ( .B1(n15501), .B2(n14945), .C1(n15635), .C2(n14942), .A(
        n2682), .ZN(n2681) );
  AOI22_X1 U2290 ( .A1(n14939), .A2(n9661), .B1(n14936), .B2(n3215), .ZN(n2682) );
  OAI221_X1 U2291 ( .B1(n15500), .B2(n14945), .C1(n15634), .C2(n14942), .A(
        n2664), .ZN(n2663) );
  AOI22_X1 U2292 ( .A1(n14939), .A2(n9662), .B1(n14935), .B2(n3230), .ZN(n2664) );
  OAI221_X1 U2293 ( .B1(n15522), .B2(n14945), .C1(n15550), .C2(n14942), .A(
        n2646), .ZN(n2645) );
  AOI22_X1 U2294 ( .A1(n14939), .A2(n9603), .B1(n14935), .B2(n3710), .ZN(n2646) );
  OAI221_X1 U2295 ( .B1(n15893), .B2(n14897), .C1(n15608), .C2(n14894), .A(
        n2654), .ZN(n2653) );
  AOI22_X1 U2296 ( .A1(n14891), .A2(n3925), .B1(n14889), .B2(Data_in[28]), 
        .ZN(n2654) );
  OAI221_X1 U2297 ( .B1(n15510), .B2(n14945), .C1(n15742), .C2(n14942), .A(
        n2628), .ZN(n2627) );
  AOI22_X1 U2298 ( .A1(n14939), .A2(n3293), .B1(n14935), .B2(n3282), .ZN(n2628) );
  OAI221_X1 U2299 ( .B1(n15892), .B2(n14897), .C1(n9438), .C2(n14894), .A(
        n2636), .ZN(n2635) );
  AOI22_X1 U2300 ( .A1(n14891), .A2(n3850), .B1(n14889), .B2(Data_in[29]), 
        .ZN(n2636) );
  OAI221_X1 U2301 ( .B1(n15521), .B2(n14945), .C1(n15431), .C2(n14942), .A(
        n2610), .ZN(n2609) );
  AOI22_X1 U2302 ( .A1(n14939), .A2(n3324), .B1(n14935), .B2(n3323), .ZN(n2610) );
  OAI221_X1 U2303 ( .B1(n3346), .B2(n14884), .C1(n16166), .C2(n14881), .A(
        n2961), .ZN(n2958) );
  AOI22_X1 U2304 ( .A1(n14878), .A2(n3722), .B1(n14877), .B2(n15378), .ZN(
        n2961) );
  OAI221_X1 U2305 ( .B1(n3347), .B2(n14884), .C1(n16165), .C2(n14881), .A(
        n2943), .ZN(n2940) );
  AOI22_X1 U2306 ( .A1(n14878), .A2(n3259), .B1(n14877), .B2(n15377), .ZN(
        n2943) );
  OAI221_X1 U2307 ( .B1(n3348), .B2(n14885), .C1(n16164), .C2(n14882), .A(
        n2781), .ZN(n2778) );
  AOI22_X1 U2308 ( .A1(n14879), .A2(n3721), .B1(n14876), .B2(n15376), .ZN(
        n2781) );
  OAI221_X1 U2309 ( .B1(n16096), .B2(n14934), .C1(n15596), .C2(n14931), .A(
        n1423), .ZN(n1417) );
  AOI22_X1 U2310 ( .A1(n14928), .A2(n15490), .B1(n14923), .B2(n15425), .ZN(
        n1423) );
  OAI221_X1 U2311 ( .B1(n15891), .B2(n14886), .C1(n16147), .C2(n14883), .A(
        n1433), .ZN(n1428) );
  AOI22_X1 U2312 ( .A1(n14880), .A2(n9650), .B1(n14875), .B2(n9769), .ZN(n1433) );
  OAI221_X1 U2313 ( .B1(n15960), .B2(n14934), .C1(n15730), .C2(n14931), .A(
        n1382), .ZN(n1342) );
  AOI22_X1 U2314 ( .A1(n14928), .A2(n9421), .B1(n14923), .B2(n9803), .ZN(n1382) );
  OAI221_X1 U2315 ( .B1(n15852), .B2(n14886), .C1(n16140), .C2(n14883), .A(
        n1403), .ZN(n1395) );
  AOI22_X1 U2316 ( .A1(n14880), .A2(n3349), .B1(n14875), .B2(n9500), .ZN(n1403) );
  OAI221_X1 U2317 ( .B1(n15980), .B2(n14934), .C1(n15623), .C2(n14931), .A(
        n1316), .ZN(n1312) );
  AOI22_X1 U2318 ( .A1(n14928), .A2(n9847), .B1(n14923), .B2(n15424), .ZN(
        n1316) );
  OAI221_X1 U2319 ( .B1(n15832), .B2(n14886), .C1(n16083), .C2(n14883), .A(
        n1333), .ZN(n1324) );
  AOI22_X1 U2320 ( .A1(n14880), .A2(n3247), .B1(n14875), .B2(n9745), .ZN(n1333) );
  OAI221_X1 U2321 ( .B1(n16095), .B2(n14934), .C1(n15535), .C2(n14931), .A(
        n1296), .ZN(n1291) );
  AOI22_X1 U2322 ( .A1(n14928), .A2(n9851), .B1(n14923), .B2(n9481), .ZN(n1296) );
  OAI221_X1 U2323 ( .B1(n15831), .B2(n14886), .C1(n16082), .C2(n14883), .A(
        n1305), .ZN(n1301) );
  AOI22_X1 U2324 ( .A1(n14880), .A2(n3628), .B1(n14875), .B2(n15464), .ZN(
        n1305) );
  OAI221_X1 U2325 ( .B1(n15979), .B2(n14934), .C1(n15595), .C2(n14931), .A(
        n1275), .ZN(n1269) );
  AOI22_X1 U2326 ( .A1(n14928), .A2(n9558), .B1(n14923), .B2(n15423), .ZN(
        n1275) );
  OAI221_X1 U2327 ( .B1(n15771), .B2(n14886), .C1(n16071), .C2(n14883), .A(
        n1284), .ZN(n1280) );
  AOI22_X1 U2328 ( .A1(n14880), .A2(n3216), .B1(n14875), .B2(n9776), .ZN(n1284) );
  OAI221_X1 U2329 ( .B1(n16094), .B2(n14934), .C1(n15594), .C2(n14931), .A(
        n1229), .ZN(n1222) );
  AOI22_X1 U2330 ( .A1(n14928), .A2(n15489), .B1(n14923), .B2(n15422), .ZN(
        n1229) );
  OAI221_X1 U2331 ( .B1(n15890), .B2(n14886), .C1(n16146), .C2(n14883), .A(
        n1252), .ZN(n1239) );
  AOI22_X1 U2332 ( .A1(n14880), .A2(n9653), .B1(n14875), .B2(n9770), .ZN(n1252) );
  OAI221_X1 U2333 ( .B1(n15978), .B2(n14934), .C1(n15593), .C2(n14931), .A(
        n1141), .ZN(n1132) );
  AOI22_X1 U2334 ( .A1(n14928), .A2(n9559), .B1(n14923), .B2(n15421), .ZN(
        n1141) );
  OAI221_X1 U2335 ( .B1(n15770), .B2(n14886), .C1(n16070), .C2(n14883), .A(
        n1171), .ZN(n1158) );
  AOI22_X1 U2336 ( .A1(n14880), .A2(n3217), .B1(n14875), .B2(n9777), .ZN(n1171) );
  OAI221_X1 U2337 ( .B1(n15949), .B2(n14934), .C1(n15533), .C2(n14931), .A(
        n2593), .ZN(n2590) );
  AOI22_X1 U2338 ( .A1(n14928), .A2(n9556), .B1(n14923), .B2(n15460), .ZN(
        n2593) );
  OAI221_X1 U2339 ( .B1(n15817), .B2(n14886), .C1(n15933), .C2(n14883), .A(
        n2601), .ZN(n2598) );
  AOI22_X1 U2340 ( .A1(n14880), .A2(n3649), .B1(n14875), .B2(n9394), .ZN(n2601) );
  OAI221_X1 U2341 ( .B1(n15954), .B2(n14932), .C1(n15673), .C2(n14929), .A(
        n3030), .ZN(n3022) );
  AOI22_X1 U2342 ( .A1(n14926), .A2(n9852), .B1(n14925), .B2(n9482), .ZN(n3030) );
  OAI221_X1 U2343 ( .B1(n15830), .B2(n14884), .C1(n15936), .C2(n14881), .A(
        n3045), .ZN(n3042) );
  AOI22_X1 U2344 ( .A1(n14878), .A2(n3944), .B1(n14877), .B2(n15379), .ZN(
        n3045) );
  OAI221_X1 U2345 ( .B1(n15953), .B2(n14932), .C1(n15672), .C2(n14929), .A(
        n3007), .ZN(n3004) );
  AOI22_X1 U2346 ( .A1(n14926), .A2(n9853), .B1(n14925), .B2(n9483), .ZN(n3007) );
  OAI221_X1 U2347 ( .B1(n15829), .B2(n14884), .C1(n15935), .C2(n14881), .A(
        n3015), .ZN(n3012) );
  AOI22_X1 U2348 ( .A1(n14878), .A2(n9683), .B1(n14877), .B2(n15462), .ZN(
        n3015) );
  OAI221_X1 U2349 ( .B1(n16038), .B2(n14932), .C1(n15671), .C2(n14929), .A(
        n2989), .ZN(n2986) );
  AOI22_X1 U2350 ( .A1(n14926), .A2(n15481), .B1(n14925), .B2(n15420), .ZN(
        n2989) );
  OAI221_X1 U2351 ( .B1(n15769), .B2(n14884), .C1(n16069), .C2(n14881), .A(
        n2997), .ZN(n2994) );
  AOI22_X1 U2352 ( .A1(n14878), .A2(n3220), .B1(n14877), .B2(n9778), .ZN(n2997) );
  OAI221_X1 U2353 ( .B1(n15977), .B2(n14932), .C1(n15622), .C2(n14929), .A(
        n2971), .ZN(n2968) );
  AOI22_X1 U2354 ( .A1(n14926), .A2(n9848), .B1(n14925), .B2(n15419), .ZN(
        n2971) );
  OAI221_X1 U2355 ( .B1(n15828), .B2(n14884), .C1(n16081), .C2(n14881), .A(
        n2979), .ZN(n2976) );
  AOI22_X1 U2356 ( .A1(n14878), .A2(n3248), .B1(n14877), .B2(n9751), .ZN(n2979) );
  OAI221_X1 U2357 ( .B1(n16127), .B2(n14932), .C1(n9721), .C2(n14929), .A(
        n2953), .ZN(n2950) );
  AOI22_X1 U2358 ( .A1(n14926), .A2(n15494), .B1(n14925), .B2(n15418), .ZN(
        n2953) );
  OAI221_X1 U2359 ( .B1(n16126), .B2(n14932), .C1(n9722), .C2(n14929), .A(
        n2935), .ZN(n2932) );
  AOI22_X1 U2360 ( .A1(n14926), .A2(n15493), .B1(n14925), .B2(n15417), .ZN(
        n2935) );
  OAI221_X1 U2361 ( .B1(n16037), .B2(n14932), .C1(n15729), .C2(n14929), .A(
        n2917), .ZN(n2914) );
  AOI22_X1 U2362 ( .A1(n14926), .A2(n15492), .B1(n14925), .B2(n15452), .ZN(
        n2917) );
  OAI221_X1 U2363 ( .B1(n15851), .B2(n14884), .C1(n15922), .C2(n14881), .A(
        n2925), .ZN(n2922) );
  AOI22_X1 U2364 ( .A1(n14878), .A2(n3265), .B1(n14877), .B2(n9336), .ZN(n2925) );
  OAI221_X1 U2365 ( .B1(n15931), .B2(n14932), .C1(n15560), .C2(n14929), .A(
        n2899), .ZN(n2896) );
  AOI22_X1 U2366 ( .A1(n14926), .A2(n15480), .B1(n14925), .B2(n9754), .ZN(
        n2899) );
  OAI221_X1 U2367 ( .B1(n15768), .B2(n14884), .C1(n16068), .C2(n14881), .A(
        n2907), .ZN(n2904) );
  AOI22_X1 U2368 ( .A1(n14878), .A2(n3218), .B1(n14877), .B2(n9779), .ZN(n2907) );
  OAI221_X1 U2369 ( .B1(n16048), .B2(n14932), .C1(n15728), .C2(n14929), .A(
        n2881), .ZN(n2878) );
  AOI22_X1 U2370 ( .A1(n14926), .A2(n9418), .B1(n14924), .B2(n9741), .ZN(n2881) );
  OAI221_X1 U2371 ( .B1(n15827), .B2(n14884), .C1(n16080), .C2(n14881), .A(
        n2889), .ZN(n2886) );
  AOI22_X1 U2372 ( .A1(n14878), .A2(n3249), .B1(n14876), .B2(n9746), .ZN(n2889) );
  OAI221_X1 U2373 ( .B1(n15910), .B2(n14884), .C1(n16032), .C2(n14881), .A(
        n2871), .ZN(n2868) );
  AOI22_X1 U2374 ( .A1(n14878), .A2(n3262), .B1(n14876), .B2(n9363), .ZN(n2871) );
  OAI221_X1 U2375 ( .B1(n15976), .B2(n14932), .C1(n15592), .C2(n14929), .A(
        n2845), .ZN(n2842) );
  AOI22_X1 U2376 ( .A1(n14926), .A2(n9560), .B1(n14924), .B2(n15415), .ZN(
        n2845) );
  OAI221_X1 U2377 ( .B1(n15909), .B2(n14884), .C1(n16145), .C2(n14881), .A(
        n2853), .ZN(n2850) );
  AOI22_X1 U2378 ( .A1(n14878), .A2(n3263), .B1(n14876), .B2(n9759), .ZN(n2853) );
  OAI221_X1 U2379 ( .B1(n16093), .B2(n14932), .C1(n15591), .C2(n14929), .A(
        n2827), .ZN(n2824) );
  AOI22_X1 U2380 ( .A1(n14926), .A2(n15487), .B1(n14924), .B2(n15414), .ZN(
        n2827) );
  OAI221_X1 U2381 ( .B1(n15889), .B2(n14884), .C1(n16144), .C2(n14881), .A(
        n2835), .ZN(n2832) );
  AOI22_X1 U2382 ( .A1(n14878), .A2(n9652), .B1(n14876), .B2(n9771), .ZN(n2835) );
  OAI221_X1 U2383 ( .B1(n16047), .B2(n14933), .C1(n15727), .C2(n14930), .A(
        n2809), .ZN(n2806) );
  AOI22_X1 U2384 ( .A1(n14927), .A2(n9419), .B1(n14924), .B2(n9742), .ZN(n2809) );
  OAI221_X1 U2385 ( .B1(n15826), .B2(n14885), .C1(n16079), .C2(n14882), .A(
        n2817), .ZN(n2814) );
  AOI22_X1 U2386 ( .A1(n14879), .A2(n3250), .B1(n14876), .B2(n9747), .ZN(n2817) );
  OAI221_X1 U2387 ( .B1(n15961), .B2(n14933), .C1(n15638), .C2(n14930), .A(
        n2791), .ZN(n2788) );
  AOI22_X1 U2388 ( .A1(n14927), .A2(n15479), .B1(n14924), .B2(n9765), .ZN(
        n2791) );
  OAI221_X1 U2389 ( .B1(n15905), .B2(n14885), .C1(n16067), .C2(n14882), .A(
        n2799), .ZN(n2796) );
  AOI22_X1 U2390 ( .A1(n14879), .A2(n3723), .B1(n14876), .B2(n9524), .ZN(n2799) );
  OAI221_X1 U2391 ( .B1(n16125), .B2(n14933), .C1(n9723), .C2(n14930), .A(
        n2773), .ZN(n2770) );
  AOI22_X1 U2392 ( .A1(n14927), .A2(n15491), .B1(n14924), .B2(n15413), .ZN(
        n2773) );
  OAI221_X1 U2393 ( .B1(n16092), .B2(n14933), .C1(n15590), .C2(n14930), .A(
        n2755), .ZN(n2752) );
  AOI22_X1 U2394 ( .A1(n14927), .A2(n15486), .B1(n14924), .B2(n15412), .ZN(
        n2755) );
  OAI221_X1 U2395 ( .B1(n15888), .B2(n14885), .C1(n16143), .C2(n14882), .A(
        n2763), .ZN(n2760) );
  AOI22_X1 U2396 ( .A1(n14879), .A2(n9648), .B1(n14876), .B2(n9772), .ZN(n2763) );
  OAI221_X1 U2397 ( .B1(n15908), .B2(n14885), .C1(n16031), .C2(n14882), .A(
        n2745), .ZN(n2742) );
  AOI22_X1 U2398 ( .A1(n14879), .A2(n3679), .B1(n14876), .B2(n9362), .ZN(n2745) );
  OAI221_X1 U2399 ( .B1(n16091), .B2(n14933), .C1(n15589), .C2(n14930), .A(
        n2719), .ZN(n2716) );
  AOI22_X1 U2400 ( .A1(n14927), .A2(n15484), .B1(n14924), .B2(n15410), .ZN(
        n2719) );
  OAI221_X1 U2401 ( .B1(n15887), .B2(n14885), .C1(n16142), .C2(n14882), .A(
        n2727), .ZN(n2724) );
  AOI22_X1 U2402 ( .A1(n14879), .A2(n9651), .B1(n14876), .B2(n9773), .ZN(n2727) );
  OAI221_X1 U2403 ( .B1(n16046), .B2(n14933), .C1(n15726), .C2(n14930), .A(
        n2701), .ZN(n2698) );
  AOI22_X1 U2404 ( .A1(n14927), .A2(n9420), .B1(n14924), .B2(n9743), .ZN(n2701) );
  OAI221_X1 U2405 ( .B1(n15825), .B2(n14885), .C1(n16078), .C2(n14882), .A(
        n2709), .ZN(n2706) );
  AOI22_X1 U2406 ( .A1(n14879), .A2(n3251), .B1(n14876), .B2(n9749), .ZN(n2709) );
  OAI221_X1 U2407 ( .B1(n15975), .B2(n14933), .C1(n15621), .C2(n14930), .A(
        n2683), .ZN(n2680) );
  AOI22_X1 U2408 ( .A1(n14927), .A2(n9849), .B1(n14924), .B2(n15409), .ZN(
        n2683) );
  OAI221_X1 U2409 ( .B1(n15824), .B2(n14885), .C1(n16077), .C2(n14882), .A(
        n2691), .ZN(n2688) );
  AOI22_X1 U2410 ( .A1(n14879), .A2(n3252), .B1(n14876), .B2(n9748), .ZN(n2691) );
  OAI221_X1 U2411 ( .B1(n15974), .B2(n14933), .C1(n15620), .C2(n14930), .A(
        n2665), .ZN(n2662) );
  AOI22_X1 U2412 ( .A1(n14927), .A2(n9850), .B1(n14923), .B2(n15408), .ZN(
        n2665) );
  OAI221_X1 U2413 ( .B1(n15823), .B2(n14885), .C1(n16076), .C2(n14882), .A(
        n2673), .ZN(n2670) );
  AOI22_X1 U2414 ( .A1(n14879), .A2(n3253), .B1(n14875), .B2(n9750), .ZN(n2673) );
  OAI221_X1 U2415 ( .B1(n16090), .B2(n14933), .C1(n15588), .C2(n14930), .A(
        n2647), .ZN(n2644) );
  AOI22_X1 U2416 ( .A1(n14927), .A2(n15483), .B1(n14923), .B2(n15407), .ZN(
        n2647) );
  OAI221_X1 U2417 ( .B1(n15886), .B2(n14885), .C1(n16141), .C2(n14882), .A(
        n2655), .ZN(n2652) );
  AOI22_X1 U2418 ( .A1(n14879), .A2(n9649), .B1(n14875), .B2(n9774), .ZN(n2655) );
  OAI221_X1 U2419 ( .B1(n16124), .B2(n14933), .C1(n15564), .C2(n14930), .A(
        n2629), .ZN(n2626) );
  AOI22_X1 U2420 ( .A1(n14927), .A2(n9873), .B1(n14923), .B2(n9498), .ZN(n2629) );
  OAI221_X1 U2421 ( .B1(n15850), .B2(n14885), .C1(n16139), .C2(n14882), .A(
        n2637), .ZN(n2634) );
  AOI22_X1 U2422 ( .A1(n14879), .A2(n3266), .B1(n14875), .B2(n9775), .ZN(n2637) );
  OAI221_X1 U2423 ( .B1(n15950), .B2(n14933), .C1(n15534), .C2(n14930), .A(
        n2611), .ZN(n2608) );
  AOI22_X1 U2424 ( .A1(n14927), .A2(n9555), .B1(n14923), .B2(n15461), .ZN(
        n2611) );
  OAI221_X1 U2425 ( .B1(n15818), .B2(n14885), .C1(n15934), .C2(n14882), .A(
        n2619), .ZN(n2616) );
  AOI22_X1 U2426 ( .A1(n14879), .A2(n3873), .B1(n14875), .B2(n9393), .ZN(n2619) );
  OAI221_X1 U2427 ( .B1(n3979), .B2(n14872), .C1(n15951), .C2(n14869), .A(
        n3016), .ZN(n3011) );
  AOI22_X1 U2428 ( .A1(n14866), .A2(n3241), .B1(n14865), .B2(n15403), .ZN(
        n3016) );
  OAI221_X1 U2429 ( .B1(n15948), .B2(n14922), .C1(n15630), .C2(n14919), .A(
        n1424), .ZN(n1416) );
  AOI22_X1 U2430 ( .A1(n14916), .A2(n15367), .B1(n14911), .B2(n15361), .ZN(
        n1424) );
  OAI221_X1 U2431 ( .B1(n16290), .B2(n14874), .C1(n16138), .C2(n14871), .A(
        n1434), .ZN(n1427) );
  AOI22_X1 U2432 ( .A1(n14868), .A2(n3236), .B1(n14863), .B2(n9841), .ZN(n1434) );
  OAI221_X1 U2433 ( .B1(n15921), .B2(n14922), .C1(n15747), .C2(n14919), .A(
        n1384), .ZN(n1341) );
  AOI22_X1 U2434 ( .A1(n14916), .A2(n9881), .B1(n14911), .B2(n15360), .ZN(
        n1384) );
  OAI221_X1 U2435 ( .B1(n16207), .B2(n14874), .C1(n15955), .C2(n14871), .A(
        n1410), .ZN(n1393) );
  AOI22_X1 U2436 ( .A1(n14868), .A2(n3237), .B1(n14863), .B2(n9863), .ZN(n1410) );
  OAI221_X1 U2437 ( .B1(n16023), .B2(n14922), .C1(n15558), .C2(n14919), .A(
        n1317), .ZN(n1311) );
  AOI22_X1 U2438 ( .A1(n14916), .A2(n9548), .B1(n14911), .B2(n9366), .ZN(n1317) );
  OAI221_X1 U2439 ( .B1(n16227), .B2(n14874), .C1(n15930), .C2(n14871), .A(
        n1334), .ZN(n1322) );
  AOI22_X1 U2440 ( .A1(n14868), .A2(n3211), .B1(n14863), .B2(n15406), .ZN(
        n1334) );
  OAI221_X1 U2441 ( .B1(n16022), .B2(n14922), .C1(n15753), .C2(n14919), .A(
        n1297), .ZN(n1290) );
  AOI22_X1 U2442 ( .A1(n14916), .A2(n9882), .B1(n14911), .B2(n9496), .ZN(n1297) );
  OAI221_X1 U2443 ( .B1(n16226), .B2(n14874), .C1(n16123), .C2(n14871), .A(
        n1306), .ZN(n1300) );
  AOI22_X1 U2444 ( .A1(n14868), .A2(n3238), .B1(n14863), .B2(n15451), .ZN(
        n1306) );
  OAI221_X1 U2445 ( .B1(n15947), .B2(n14922), .C1(n15741), .C2(n14919), .A(
        n1276), .ZN(n1268) );
  AOI22_X1 U2446 ( .A1(n14916), .A2(n9876), .B1(n14911), .B2(n9396), .ZN(n1276) );
  OAI221_X1 U2447 ( .B1(n16252), .B2(n14874), .C1(n16030), .C2(n14871), .A(
        n1285), .ZN(n1279) );
  AOI22_X1 U2448 ( .A1(n14868), .A2(n3219), .B1(n14863), .B2(n15405), .ZN(
        n1285) );
  OAI221_X1 U2449 ( .B1(n15946), .B2(n14922), .C1(n15629), .C2(n14919), .A(
        n1230), .ZN(n1213) );
  AOI22_X1 U2450 ( .A1(n14916), .A2(n15366), .B1(n14911), .B2(n15359), .ZN(
        n1230) );
  OAI221_X1 U2451 ( .B1(n16289), .B2(n14874), .C1(n16137), .C2(n14871), .A(
        n1255), .ZN(n1234) );
  AOI22_X1 U2452 ( .A1(n14868), .A2(n3239), .B1(n14863), .B2(n9842), .ZN(n1255) );
  OAI221_X1 U2453 ( .B1(n15945), .B2(n14922), .C1(n15740), .C2(n14919), .A(
        n1146), .ZN(n1131) );
  AOI22_X1 U2454 ( .A1(n14916), .A2(n9877), .B1(n14911), .B2(n9399), .ZN(n1146) );
  OAI221_X1 U2455 ( .B1(n16251), .B2(n14874), .C1(n16029), .C2(n14871), .A(
        n1182), .ZN(n1157) );
  AOI22_X1 U2456 ( .A1(n14868), .A2(n3264), .B1(n14863), .B2(n15404), .ZN(
        n1182) );
  OAI221_X1 U2457 ( .B1(n15923), .B2(n14922), .C1(n15561), .C2(n14919), .A(
        n2594), .ZN(n2589) );
  AOI22_X1 U2458 ( .A1(n14916), .A2(n9880), .B1(n14911), .B2(n9365), .ZN(n2594) );
  OAI221_X1 U2459 ( .B1(n16283), .B2(n14874), .C1(n16033), .C2(n14871), .A(
        n2602), .ZN(n2597) );
  AOI22_X1 U2460 ( .A1(n14868), .A2(n9685), .B1(n14863), .B2(n15453), .ZN(
        n2602) );
  OAI221_X1 U2461 ( .B1(n9597), .B2(n14910), .C1(n15713), .C2(n14907), .A(
        n1425), .ZN(n1415) );
  AOI22_X1 U2462 ( .A1(n14904), .A2(n9671), .B1(n14899), .B2(n3117), .ZN(n1425) );
  OAI221_X1 U2463 ( .B1(n9596), .B2(n14910), .C1(n15711), .C2(n14907), .A(
        n1231), .ZN(n1212) );
  AOI22_X1 U2464 ( .A1(n14904), .A2(n9669), .B1(n14899), .B2(n3118), .ZN(n1231) );
  OAI221_X1 U2465 ( .B1(n3629), .B2(n14908), .C1(n9574), .C2(n14905), .A(n2955), .ZN(n2948) );
  AOI22_X1 U2466 ( .A1(n14902), .A2(n3976), .B1(n14901), .B2(n15467), .ZN(
        n2955) );
  OAI221_X1 U2467 ( .B1(n3630), .B2(n14908), .C1(n9573), .C2(n14905), .A(n2937), .ZN(n2930) );
  AOI22_X1 U2468 ( .A1(n14902), .A2(n3977), .B1(n14901), .B2(n15466), .ZN(
        n2937) );
  OAI221_X1 U2469 ( .B1(n9593), .B2(n14908), .C1(n15706), .C2(n14905), .A(
        n2829), .ZN(n2822) );
  AOI22_X1 U2470 ( .A1(n14902), .A2(n9667), .B1(n14900), .B2(n3119), .ZN(n2829) );
  OAI221_X1 U2471 ( .B1(n9439), .B2(n14909), .C1(n15833), .C2(n14906), .A(
        n2793), .ZN(n2786) );
  AOI22_X1 U2472 ( .A1(n14903), .A2(n3053), .B1(n14900), .B2(n3091), .ZN(n2793) );
  OAI221_X1 U2473 ( .B1(n3631), .B2(n14909), .C1(n9575), .C2(n14906), .A(n2775), .ZN(n2768) );
  AOI22_X1 U2474 ( .A1(n14903), .A2(n3978), .B1(n14900), .B2(n15465), .ZN(
        n2775) );
  OAI221_X1 U2475 ( .B1(n9595), .B2(n14909), .C1(n15705), .C2(n14906), .A(
        n2757), .ZN(n2750) );
  AOI22_X1 U2476 ( .A1(n14903), .A2(n9668), .B1(n14900), .B2(n3120), .ZN(n2757) );
  OAI221_X1 U2477 ( .B1(n9594), .B2(n14909), .C1(n15704), .C2(n14906), .A(
        n2721), .ZN(n2714) );
  AOI22_X1 U2478 ( .A1(n14903), .A2(n9673), .B1(n14900), .B2(n3121), .ZN(n2721) );
  OAI221_X1 U2479 ( .B1(n9451), .B2(n14909), .C1(n15703), .C2(n14906), .A(
        n2649), .ZN(n2642) );
  AOI22_X1 U2480 ( .A1(n14903), .A2(n9672), .B1(n14899), .B2(n3122), .ZN(n2649) );
  OAI221_X1 U2481 ( .B1(n15667), .B2(n14910), .C1(n15775), .C2(n14907), .A(
        n1387), .ZN(n1340) );
  AOI22_X1 U2482 ( .A1(n14904), .A2(n3124), .B1(n14899), .B2(n3962), .ZN(n1387) );
  OAI221_X1 U2483 ( .B1(n15666), .B2(n14910), .C1(n15779), .C2(n14907), .A(
        n1319), .ZN(n1310) );
  AOI22_X1 U2484 ( .A1(n14904), .A2(n3167), .B1(n14899), .B2(n3125), .ZN(n1319) );
  OAI221_X1 U2485 ( .B1(n15665), .B2(n14910), .C1(n15767), .C2(n14907), .A(
        n1298), .ZN(n1289) );
  AOI22_X1 U2486 ( .A1(n14904), .A2(n3970), .B1(n14899), .B2(n3126), .ZN(n1298) );
  OAI221_X1 U2487 ( .B1(n15696), .B2(n14910), .C1(n15712), .C2(n14907), .A(
        n1277), .ZN(n1265) );
  AOI22_X1 U2488 ( .A1(n14904), .A2(n3132), .B1(n14899), .B2(n3713), .ZN(n1277) );
  OAI221_X1 U2489 ( .B1(n15695), .B2(n14910), .C1(n15710), .C2(n14907), .A(
        n1151), .ZN(n1130) );
  AOI22_X1 U2490 ( .A1(n14904), .A2(n3133), .B1(n14899), .B2(n3704), .ZN(n1151) );
  OAI221_X1 U2491 ( .B1(n15843), .B2(n14910), .C1(n15754), .C2(n14907), .A(
        n2595), .ZN(n2588) );
  AOI22_X1 U2492 ( .A1(n14904), .A2(n3134), .B1(n14899), .B2(n3149), .ZN(n2595) );
  OAI221_X1 U2493 ( .B1(n15926), .B2(n14920), .C1(n15543), .C2(n14917), .A(
        n3035), .ZN(n3021) );
  AOI22_X1 U2494 ( .A1(n14914), .A2(n9862), .B1(n14913), .B2(n9470), .ZN(n3035) );
  OAI221_X1 U2495 ( .B1(n16306), .B2(n14872), .C1(n15952), .C2(n14869), .A(
        n3046), .ZN(n3041) );
  AOI22_X1 U2496 ( .A1(n14866), .A2(n3321), .B1(n14865), .B2(n15478), .ZN(
        n3046) );
  OAI221_X1 U2497 ( .B1(n15925), .B2(n14920), .C1(n15597), .C2(n14917), .A(
        n3008), .ZN(n3003) );
  AOI22_X1 U2498 ( .A1(n14914), .A2(n9883), .B1(n14913), .B2(n9497), .ZN(n3008) );
  OAI221_X1 U2499 ( .B1(n15944), .B2(n14920), .C1(n15739), .C2(n14917), .A(
        n2990), .ZN(n2985) );
  AOI22_X1 U2500 ( .A1(n14914), .A2(n9866), .B1(n14913), .B2(n9397), .ZN(n2990) );
  OAI221_X1 U2501 ( .B1(n16250), .B2(n14872), .C1(n16028), .C2(n14869), .A(
        n2998), .ZN(n2993) );
  AOI22_X1 U2502 ( .A1(n14866), .A2(n3268), .B1(n14865), .B2(n9864), .ZN(n2998) );
  OAI221_X1 U2503 ( .B1(n16021), .B2(n14920), .C1(n15644), .C2(n14917), .A(
        n2972), .ZN(n2967) );
  AOI22_X1 U2504 ( .A1(n14914), .A2(n9552), .B1(n14913), .B2(n9371), .ZN(n2972) );
  OAI221_X1 U2505 ( .B1(n16225), .B2(n14872), .C1(n15929), .C2(n14869), .A(
        n2980), .ZN(n2975) );
  AOI22_X1 U2506 ( .A1(n14866), .A2(n3276), .B1(n14865), .B2(n15402), .ZN(
        n2980) );
  OAI221_X1 U2507 ( .B1(n16066), .B2(n14920), .C1(n15437), .C2(n14917), .A(
        n2954), .ZN(n2949) );
  AOI22_X1 U2508 ( .A1(n14914), .A2(n15477), .B1(n14913), .B2(n15473), .ZN(
        n2954) );
  OAI221_X1 U2509 ( .B1(n16313), .B2(n14872), .C1(n16075), .C2(n14869), .A(
        n2962), .ZN(n2957) );
  AOI22_X1 U2510 ( .A1(n14866), .A2(n3277), .B1(n14865), .B2(n15401), .ZN(
        n2962) );
  OAI221_X1 U2511 ( .B1(n16065), .B2(n14920), .C1(n15436), .C2(n14917), .A(
        n2936), .ZN(n2931) );
  AOI22_X1 U2512 ( .A1(n14914), .A2(n15476), .B1(n14913), .B2(n15472), .ZN(
        n2936) );
  OAI221_X1 U2513 ( .B1(n16312), .B2(n14872), .C1(n16074), .C2(n14869), .A(
        n2944), .ZN(n2939) );
  AOI22_X1 U2514 ( .A1(n14866), .A2(n3278), .B1(n14865), .B2(n15400), .ZN(
        n2944) );
  OAI221_X1 U2515 ( .B1(n16163), .B2(n14920), .C1(n15746), .C2(n14917), .A(
        n2918), .ZN(n2913) );
  AOI22_X1 U2516 ( .A1(n14914), .A2(n9826), .B1(n14913), .B2(n9401), .ZN(n2918) );
  OAI221_X1 U2517 ( .B1(n16206), .B2(n14872), .C1(n15932), .C2(n14869), .A(
        n2926), .ZN(n2921) );
  AOI22_X1 U2518 ( .A1(n14866), .A2(n3280), .B1(n14865), .B2(n9562), .ZN(n2926) );
  OAI221_X1 U2519 ( .B1(n15943), .B2(n14920), .C1(n15738), .C2(n14917), .A(
        n2900), .ZN(n2895) );
  AOI22_X1 U2520 ( .A1(n14914), .A2(n9878), .B1(n14913), .B2(n9400), .ZN(n2900) );
  OAI221_X1 U2521 ( .B1(n16249), .B2(n14872), .C1(n16027), .C2(n14869), .A(
        n2908), .ZN(n2903) );
  AOI22_X1 U2522 ( .A1(n14866), .A2(n3275), .B1(n14865), .B2(n15450), .ZN(
        n2908) );
  OAI221_X1 U2523 ( .B1(n16020), .B2(n14920), .C1(n15643), .C2(n14917), .A(
        n2882), .ZN(n2877) );
  AOI22_X1 U2524 ( .A1(n14914), .A2(n9549), .B1(n14912), .B2(n9370), .ZN(n2882) );
  OAI221_X1 U2525 ( .B1(n16224), .B2(n14872), .C1(n16122), .C2(n14869), .A(
        n2890), .ZN(n2885) );
  AOI22_X1 U2526 ( .A1(n14866), .A2(n3281), .B1(n14864), .B2(n15399), .ZN(
        n2890) );
  OAI221_X1 U2527 ( .B1(n16064), .B2(n14920), .C1(n15540), .C2(n14917), .A(
        n2864), .ZN(n2859) );
  AOI22_X1 U2528 ( .A1(n14914), .A2(n9856), .B1(n14912), .B2(n9402), .ZN(n2864) );
  OAI221_X1 U2529 ( .B1(n16248), .B2(n14872), .C1(n16026), .C2(n14869), .A(
        n2872), .ZN(n2867) );
  AOI22_X1 U2530 ( .A1(n14866), .A2(n3288), .B1(n14864), .B2(n15469), .ZN(
        n2872) );
  OAI221_X1 U2531 ( .B1(n15942), .B2(n14920), .C1(n15628), .C2(n14917), .A(
        n2846), .ZN(n2841) );
  AOI22_X1 U2532 ( .A1(n14914), .A2(n9411), .B1(n14912), .B2(n9768), .ZN(n2846) );
  OAI221_X1 U2533 ( .B1(n16263), .B2(n14872), .C1(n16136), .C2(n14869), .A(
        n2854), .ZN(n2849) );
  AOI22_X1 U2534 ( .A1(n14866), .A2(n9681), .B1(n14864), .B2(n15398), .ZN(
        n2854) );
  OAI221_X1 U2535 ( .B1(n15941), .B2(n14920), .C1(n15627), .C2(n14917), .A(
        n2828), .ZN(n2823) );
  AOI22_X1 U2536 ( .A1(n14914), .A2(n15365), .B1(n14912), .B2(n15358), .ZN(
        n2828) );
  OAI221_X1 U2537 ( .B1(n16288), .B2(n14872), .C1(n16135), .C2(n14869), .A(
        n2836), .ZN(n2831) );
  AOI22_X1 U2538 ( .A1(n14866), .A2(n3243), .B1(n14864), .B2(n9843), .ZN(n2836) );
  OAI221_X1 U2539 ( .B1(n16019), .B2(n14921), .C1(n15642), .C2(n14918), .A(
        n2810), .ZN(n2805) );
  AOI22_X1 U2540 ( .A1(n14915), .A2(n9550), .B1(n14912), .B2(n9368), .ZN(n2810) );
  OAI221_X1 U2541 ( .B1(n16223), .B2(n14873), .C1(n16121), .C2(n14870), .A(
        n2818), .ZN(n2813) );
  AOI22_X1 U2542 ( .A1(n14867), .A2(n3306), .B1(n14864), .B2(n15397), .ZN(
        n2818) );
  OAI221_X1 U2543 ( .B1(n16063), .B2(n14921), .C1(n15780), .C2(n14918), .A(
        n2792), .ZN(n2787) );
  AOI22_X1 U2544 ( .A1(n14915), .A2(n15475), .B1(n14912), .B2(n15471), .ZN(
        n2792) );
  OAI221_X1 U2545 ( .B1(n16199), .B2(n14873), .C1(n16025), .C2(n14870), .A(
        n2800), .ZN(n2795) );
  AOI22_X1 U2546 ( .A1(n14867), .A2(n3307), .B1(n14864), .B2(n9874), .ZN(n2800) );
  OAI221_X1 U2547 ( .B1(n16062), .B2(n14921), .C1(n15435), .C2(n14918), .A(
        n2774), .ZN(n2769) );
  AOI22_X1 U2548 ( .A1(n14915), .A2(n15474), .B1(n14912), .B2(n15470), .ZN(
        n2774) );
  OAI221_X1 U2549 ( .B1(n16311), .B2(n14873), .C1(n16073), .C2(n14870), .A(
        n2782), .ZN(n2777) );
  AOI22_X1 U2550 ( .A1(n14867), .A2(n3309), .B1(n14864), .B2(n15396), .ZN(
        n2782) );
  OAI221_X1 U2551 ( .B1(n15940), .B2(n14921), .C1(n15626), .C2(n14918), .A(
        n2756), .ZN(n2751) );
  AOI22_X1 U2552 ( .A1(n14915), .A2(n15364), .B1(n14912), .B2(n15357), .ZN(
        n2756) );
  OAI221_X1 U2553 ( .B1(n16287), .B2(n14873), .C1(n16134), .C2(n14870), .A(
        n2764), .ZN(n2759) );
  AOI22_X1 U2554 ( .A1(n14867), .A2(n3244), .B1(n14864), .B2(n9845), .ZN(n2764) );
  OAI221_X1 U2555 ( .B1(n16061), .B2(n14921), .C1(n15539), .C2(n14918), .A(
        n2738), .ZN(n2733) );
  AOI22_X1 U2556 ( .A1(n14915), .A2(n9857), .B1(n14912), .B2(n9398), .ZN(n2738) );
  OAI221_X1 U2557 ( .B1(n16247), .B2(n14873), .C1(n16024), .C2(n14870), .A(
        n2746), .ZN(n2741) );
  AOI22_X1 U2558 ( .A1(n14867), .A2(n3315), .B1(n14864), .B2(n15468), .ZN(
        n2746) );
  OAI221_X1 U2559 ( .B1(n15939), .B2(n14921), .C1(n15625), .C2(n14918), .A(
        n2720), .ZN(n2715) );
  AOI22_X1 U2560 ( .A1(n14915), .A2(n15363), .B1(n14912), .B2(n15356), .ZN(
        n2720) );
  OAI221_X1 U2561 ( .B1(n16286), .B2(n14873), .C1(n16133), .C2(n14870), .A(
        n2728), .ZN(n2723) );
  AOI22_X1 U2562 ( .A1(n14867), .A2(n3258), .B1(n14864), .B2(n9844), .ZN(n2728) );
  OAI221_X1 U2563 ( .B1(n16018), .B2(n14921), .C1(n15641), .C2(n14918), .A(
        n2702), .ZN(n2697) );
  AOI22_X1 U2564 ( .A1(n14915), .A2(n9553), .B1(n14912), .B2(n9369), .ZN(n2702) );
  OAI221_X1 U2565 ( .B1(n16222), .B2(n14873), .C1(n16120), .C2(n14870), .A(
        n2710), .ZN(n2705) );
  AOI22_X1 U2566 ( .A1(n14867), .A2(n3317), .B1(n14864), .B2(n15395), .ZN(
        n2710) );
  OAI221_X1 U2567 ( .B1(n16017), .B2(n14921), .C1(n15640), .C2(n14918), .A(
        n2684), .ZN(n2679) );
  AOI22_X1 U2568 ( .A1(n14915), .A2(n9551), .B1(n14912), .B2(n9372), .ZN(n2684) );
  OAI221_X1 U2569 ( .B1(n16221), .B2(n14873), .C1(n15928), .C2(n14870), .A(
        n2692), .ZN(n2687) );
  AOI22_X1 U2570 ( .A1(n14867), .A2(n3319), .B1(n14864), .B2(n15394), .ZN(
        n2692) );
  OAI221_X1 U2571 ( .B1(n16016), .B2(n14921), .C1(n15639), .C2(n14918), .A(
        n2666), .ZN(n2661) );
  AOI22_X1 U2572 ( .A1(n14915), .A2(n9554), .B1(n14911), .B2(n9367), .ZN(n2666) );
  OAI221_X1 U2573 ( .B1(n16220), .B2(n14873), .C1(n15927), .C2(n14870), .A(
        n2674), .ZN(n2669) );
  AOI22_X1 U2574 ( .A1(n14867), .A2(n3331), .B1(n14863), .B2(n15393), .ZN(
        n2674) );
  OAI221_X1 U2575 ( .B1(n15938), .B2(n14921), .C1(n15624), .C2(n14918), .A(
        n2648), .ZN(n2643) );
  AOI22_X1 U2576 ( .A1(n14915), .A2(n15362), .B1(n14911), .B2(n15355), .ZN(
        n2648) );
  OAI221_X1 U2577 ( .B1(n16285), .B2(n14873), .C1(n16132), .C2(n14870), .A(
        n2656), .ZN(n2651) );
  AOI22_X1 U2578 ( .A1(n14867), .A2(n3245), .B1(n14863), .B2(n9846), .ZN(n2656) );
  OAI221_X1 U2579 ( .B1(n15937), .B2(n14921), .C1(n15559), .C2(n14918), .A(
        n2630), .ZN(n2625) );
  AOI22_X1 U2580 ( .A1(n14915), .A2(n9547), .B1(n14911), .B2(n15354), .ZN(
        n2630) );
  OAI221_X1 U2581 ( .B1(n16262), .B2(n14873), .C1(n16072), .C2(n14870), .A(
        n2638), .ZN(n2633) );
  AOI22_X1 U2582 ( .A1(n14867), .A2(n3246), .B1(n14863), .B2(n9858), .ZN(n2638) );
  OAI221_X1 U2583 ( .B1(n15924), .B2(n14921), .C1(n15562), .C2(n14918), .A(
        n2612), .ZN(n2607) );
  AOI22_X1 U2584 ( .A1(n14915), .A2(n9879), .B1(n14911), .B2(n9364), .ZN(n2612) );
  OAI221_X1 U2585 ( .B1(n16284), .B2(n14873), .C1(n16034), .C2(n14870), .A(
        n2620), .ZN(n2615) );
  AOI22_X1 U2586 ( .A1(n14867), .A2(n9684), .B1(n14863), .B2(n15454), .ZN(
        n2620) );
  OAI221_X1 U2587 ( .B1(n15863), .B2(n14908), .C1(n15766), .C2(n14905), .A(
        n3039), .ZN(n3020) );
  AOI22_X1 U2588 ( .A1(n14902), .A2(n3055), .B1(n14901), .B2(n3131), .ZN(n3039) );
  OAI221_X1 U2589 ( .B1(n15701), .B2(n14908), .C1(n15765), .C2(n14905), .A(
        n3009), .ZN(n3002) );
  AOI22_X1 U2590 ( .A1(n14902), .A2(n15445), .B1(n14901), .B2(n3150), .ZN(
        n3009) );
  OAI221_X1 U2591 ( .B1(n15806), .B2(n14908), .C1(n15709), .C2(n14905), .A(
        n2991), .ZN(n2984) );
  AOI22_X1 U2592 ( .A1(n14902), .A2(n3151), .B1(n14901), .B2(n3094), .ZN(n2991) );
  OAI221_X1 U2593 ( .B1(n15664), .B2(n14908), .C1(n15778), .C2(n14905), .A(
        n2973), .ZN(n2966) );
  AOI22_X1 U2594 ( .A1(n14902), .A2(n3152), .B1(n14901), .B2(n3168), .ZN(n2973) );
  OAI221_X1 U2595 ( .B1(n15694), .B2(n14908), .C1(n15774), .C2(n14905), .A(
        n2919), .ZN(n2912) );
  AOI22_X1 U2596 ( .A1(n14902), .A2(n3975), .B1(n14901), .B2(n3101), .ZN(n2919) );
  OAI221_X1 U2597 ( .B1(n15798), .B2(n14908), .C1(n15708), .C2(n14905), .A(
        n2901), .ZN(n2894) );
  AOI22_X1 U2598 ( .A1(n14902), .A2(n3169), .B1(n14901), .B2(n3714), .ZN(n2901) );
  OAI221_X1 U2599 ( .B1(n15663), .B2(n14908), .C1(n15764), .C2(n14905), .A(
        n2883), .ZN(n2876) );
  AOI22_X1 U2600 ( .A1(n14902), .A2(n3170), .B1(n14900), .B2(n3171), .ZN(n2883) );
  OAI221_X1 U2601 ( .B1(n15725), .B2(n14908), .C1(n15920), .C2(n14905), .A(
        n2865), .ZN(n2858) );
  AOI22_X1 U2602 ( .A1(n14902), .A2(n3972), .B1(n14900), .B2(n3650), .ZN(n2865) );
  OAI221_X1 U2603 ( .B1(n15700), .B2(n14908), .C1(n15707), .C2(n14905), .A(
        n2847), .ZN(n2840) );
  AOI22_X1 U2604 ( .A1(n14902), .A2(n3172), .B1(n14900), .B2(n3088), .ZN(n2847) );
  OAI221_X1 U2605 ( .B1(n15662), .B2(n14909), .C1(n15763), .C2(n14906), .A(
        n2811), .ZN(n2804) );
  AOI22_X1 U2606 ( .A1(n14903), .A2(n3173), .B1(n14900), .B2(n3174), .ZN(n2811) );
  OAI221_X1 U2607 ( .B1(n15724), .B2(n14909), .C1(n15919), .C2(n14906), .A(
        n2739), .ZN(n2732) );
  AOI22_X1 U2608 ( .A1(n14903), .A2(n3971), .B1(n14900), .B2(n3635), .ZN(n2739) );
  OAI221_X1 U2609 ( .B1(n15661), .B2(n14909), .C1(n15762), .C2(n14906), .A(
        n2703), .ZN(n2696) );
  AOI22_X1 U2610 ( .A1(n14903), .A2(n3176), .B1(n14900), .B2(n3177), .ZN(n2703) );
  OAI221_X1 U2611 ( .B1(n15660), .B2(n14909), .C1(n15777), .C2(n14906), .A(
        n2685), .ZN(n2678) );
  AOI22_X1 U2612 ( .A1(n14903), .A2(n3186), .B1(n14900), .B2(n3187), .ZN(n2685) );
  OAI221_X1 U2613 ( .B1(n15659), .B2(n14909), .C1(n15776), .C2(n14906), .A(
        n2667), .ZN(n2660) );
  AOI22_X1 U2614 ( .A1(n14903), .A2(n3191), .B1(n14899), .B2(n3192), .ZN(n2667) );
  OAI221_X1 U2615 ( .B1(n15699), .B2(n14909), .C1(n15702), .C2(n14906), .A(
        n2631), .ZN(n2624) );
  AOI22_X1 U2616 ( .A1(n14903), .A2(n9670), .B1(n14899), .B2(n3967), .ZN(n2631) );
  OAI221_X1 U2617 ( .B1(n15844), .B2(n14909), .C1(n15755), .C2(n14906), .A(
        n2613), .ZN(n2606) );
  AOI22_X1 U2618 ( .A1(n14903), .A2(n3196), .B1(n14899), .B2(n3148), .ZN(n2613) );
  AOI22_X1 U2619 ( .A1(n14856), .A2(n3071), .B1(n14851), .B2(n9816), .ZN(n1435) );
  AOI22_X1 U2620 ( .A1(n14856), .A2(n3078), .B1(n14851), .B2(n9817), .ZN(n1412) );
  AOI22_X1 U2621 ( .A1(n14856), .A2(n9612), .B1(n14851), .B2(n15375), .ZN(
        n1336) );
  AOI22_X1 U2622 ( .A1(n14856), .A2(n3103), .B1(n14851), .B2(n9818), .ZN(n1307) );
  AOI22_X1 U2623 ( .A1(n14856), .A2(n3057), .B1(n14851), .B2(n9813), .ZN(n1286) );
  AOI22_X1 U2624 ( .A1(n14856), .A2(n3072), .B1(n14851), .B2(n9819), .ZN(n1257) );
  AOI22_X1 U2625 ( .A1(n14856), .A2(n3058), .B1(n14851), .B2(n9814), .ZN(n1201) );
  AOI22_X1 U2626 ( .A1(n14854), .A2(n3100), .B1(n14853), .B2(n15374), .ZN(
        n3047) );
  AOI22_X1 U2627 ( .A1(n14854), .A2(n3102), .B1(n14853), .B2(n9820), .ZN(n3017) );
  AOI22_X1 U2628 ( .A1(n14854), .A2(n3059), .B1(n14853), .B2(n15459), .ZN(
        n2999) );
  AOI22_X1 U2629 ( .A1(n14854), .A2(n9613), .B1(n14853), .B2(n15373), .ZN(
        n2981) );
  AOI22_X1 U2630 ( .A1(n14854), .A2(n3128), .B1(n14853), .B2(n9867), .ZN(n2963) );
  AOI22_X1 U2631 ( .A1(n14854), .A2(n3129), .B1(n14853), .B2(n9868), .ZN(n2945) );
  AOI22_X1 U2632 ( .A1(n14854), .A2(n3099), .B1(n14853), .B2(n9854), .ZN(n2927) );
  AOI22_X1 U2633 ( .A1(n14854), .A2(n3069), .B1(n14853), .B2(n9815), .ZN(n2909) );
  AOI22_X1 U2634 ( .A1(n14854), .A2(n3105), .B1(n14852), .B2(n15372), .ZN(
        n2891) );
  AOI22_X1 U2635 ( .A1(n14854), .A2(n3108), .B1(n14852), .B2(n9870), .ZN(n2873) );
  AOI22_X1 U2636 ( .A1(n14854), .A2(n3073), .B1(n14852), .B2(n9827), .ZN(n2855) );
  AOI22_X1 U2637 ( .A1(n14854), .A2(n3074), .B1(n14852), .B2(n9821), .ZN(n2837) );
  AOI22_X1 U2638 ( .A1(n14855), .A2(n3104), .B1(n14852), .B2(n15371), .ZN(
        n2819) );
  AOI22_X1 U2639 ( .A1(n14855), .A2(n3106), .B1(n14852), .B2(n9890), .ZN(n2801) );
  AOI22_X1 U2640 ( .A1(n14855), .A2(n3130), .B1(n14852), .B2(n9869), .ZN(n2783) );
  AOI22_X1 U2641 ( .A1(n14855), .A2(n3075), .B1(n14852), .B2(n9822), .ZN(n2765) );
  AOI22_X1 U2642 ( .A1(n14855), .A2(n3109), .B1(n14852), .B2(n9871), .ZN(n2747) );
  AOI22_X1 U2643 ( .A1(n14855), .A2(n3076), .B1(n14852), .B2(n9823), .ZN(n2729) );
  AOI22_X1 U2644 ( .A1(n14855), .A2(n3107), .B1(n14852), .B2(n15370), .ZN(
        n2711) );
  AOI22_X1 U2645 ( .A1(n14855), .A2(n9614), .B1(n14852), .B2(n15369), .ZN(
        n2693) );
  AOI22_X1 U2646 ( .A1(n14855), .A2(n9615), .B1(n14851), .B2(n15368), .ZN(
        n2675) );
  AOI22_X1 U2647 ( .A1(n14855), .A2(n3077), .B1(n14851), .B2(n9824), .ZN(n2657) );
  AOI22_X1 U2648 ( .A1(n14855), .A2(n3070), .B1(n14851), .B2(n9825), .ZN(n2639) );
  AOI22_X1 U2649 ( .A1(n14855), .A2(n9656), .B1(n14851), .B2(n15458), .ZN(
        n2621) );
  AOI22_X1 U2650 ( .A1(n14856), .A2(n9655), .B1(n14851), .B2(n15457), .ZN(
        n2603) );
  INV_X1 U2651 ( .A(Read_two_address[2]), .ZN(n15282) );
  INV_X1 U2652 ( .A(Read_two_address[4]), .ZN(n15284) );
  INV_X1 U2653 ( .A(Read_two_address[3]), .ZN(n15283) );
  OAI22_X1 U2654 ( .A1(n14709), .A2(n1126), .B1(n14948), .B2(n15750), .ZN(
        n1375) );
  OAI22_X1 U2655 ( .A1(n14646), .A2(n14947), .B1(n14953), .B2(n15646), .ZN(
        n1354) );
  OAI22_X1 U2656 ( .A1(n14622), .A2(n14947), .B1(n14955), .B2(n15549), .ZN(
        n1346) );
  OAI22_X1 U2657 ( .A1(n14637), .A2(n14947), .B1(n14954), .B2(n15548), .ZN(
        n1351) );
  OAI22_X1 U2658 ( .A1(n14676), .A2(n1126), .B1(n14951), .B2(n15547), .ZN(
        n1364) );
  OAI22_X1 U2659 ( .A1(n14688), .A2(n1126), .B1(n14950), .B2(n15546), .ZN(
        n1368) );
  OAI22_X1 U2660 ( .A1(n14694), .A2(n1126), .B1(n14949), .B2(n15545), .ZN(
        n1370) );
  OAI22_X1 U2661 ( .A1(n14706), .A2(n1126), .B1(n14948), .B2(n15544), .ZN(
        n1374) );
  INV_X1 U2662 ( .A(Read_two_address[1]), .ZN(n15281) );
  INV_X1 U2663 ( .A(Read_two_address[0]), .ZN(n15280) );
  OAI22_X1 U2664 ( .A1(n15237), .A2(n16282), .B1(n1081), .B2(n14620), .ZN(
        n3482) );
  OAI22_X1 U2665 ( .A1(n15237), .A2(n16281), .B1(n1081), .B2(n14632), .ZN(
        n3480) );
  OAI22_X1 U2666 ( .A1(n15237), .A2(n16280), .B1(n1081), .B2(n14635), .ZN(
        n3479) );
  OAI22_X1 U2667 ( .A1(n15234), .A2(n16279), .B1(n1081), .B2(n14638), .ZN(
        n3624) );
  OAI22_X1 U2668 ( .A1(n15241), .A2(n16278), .B1(n14653), .B2(n15233), .ZN(
        n1293) );
  OAI22_X1 U2669 ( .A1(n15241), .A2(n16277), .B1(n14656), .B2(n1081), .ZN(
        n1294) );
  OAI22_X1 U2670 ( .A1(n15234), .A2(n16276), .B1(n1081), .B2(n14671), .ZN(
        n3623) );
  OAI22_X1 U2671 ( .A1(n15234), .A2(n16275), .B1(n1081), .B2(n14674), .ZN(
        n3622) );
  OAI22_X1 U2672 ( .A1(n15241), .A2(n16274), .B1(n14683), .B2(n1081), .ZN(
        n1303) );
  OAI22_X1 U2673 ( .A1(n15235), .A2(n16273), .B1(n1081), .B2(n14686), .ZN(
        n3621) );
  OAI22_X1 U2674 ( .A1(n15239), .A2(n16272), .B1(n1081), .B2(n14692), .ZN(
        n3474) );
  OAI22_X1 U2675 ( .A1(n15240), .A2(n16271), .B1(n1081), .B2(n14704), .ZN(
        n3470) );
  OAI22_X1 U2676 ( .A1(n15247), .A2(n16243), .B1(n15255), .B2(n14626), .ZN(
        n2052) );
  OAI22_X1 U2677 ( .A1(n15246), .A2(n16242), .B1(n15254), .B2(n14650), .ZN(
        n2060) );
  OAI22_X1 U2678 ( .A1(n15247), .A2(n16241), .B1(n15251), .B2(n14698), .ZN(
        n2076) );
  OAI22_X1 U2679 ( .A1(n15247), .A2(n16240), .B1(n15251), .B2(n14701), .ZN(
        n2077) );
  OAI22_X1 U2680 ( .A1(n15119), .A2(n16159), .B1(n14688), .B2(n15117), .ZN(
        n3577) );
  OAI22_X1 U2681 ( .A1(n15120), .A2(n16158), .B1(n14694), .B2(n15117), .ZN(
        n3576) );
  OAI22_X1 U2682 ( .A1(n15120), .A2(n16157), .B1(n14706), .B2(n15117), .ZN(
        n3575) );
  OAI22_X1 U2683 ( .A1(n15054), .A2(n16154), .B1(n14663), .B2(n15050), .ZN(
        n3504) );
  OAI22_X1 U2684 ( .A1(n15241), .A2(n16148), .B1(n1081), .B2(n14624), .ZN(
        n1283) );
  OAI22_X1 U2685 ( .A1(n15247), .A2(n16131), .B1(n15253), .B2(n14665), .ZN(
        n2065) );
  OAI22_X1 U2686 ( .A1(n15247), .A2(n16130), .B1(n15252), .B2(n14677), .ZN(
        n2069) );
  OAI22_X1 U2687 ( .A1(n15247), .A2(n16129), .B1(n15252), .B2(n14695), .ZN(
        n2075) );
  OAI22_X1 U2688 ( .A1(n15058), .A2(n16005), .B1(n14660), .B2(n15051), .ZN(
        n3389) );
  OAI22_X1 U2689 ( .A1(n15152), .A2(n15995), .B1(n15144), .B2(n14623), .ZN(
        n1635) );
  OAI22_X1 U2690 ( .A1(n15055), .A2(n15983), .B1(n14669), .B2(n15050), .ZN(
        n3502) );
  OAI22_X1 U2691 ( .A1(n15056), .A2(n15982), .B1(n14689), .B2(n15050), .ZN(
        n3499) );
  OAI22_X1 U2692 ( .A1(n15180), .A2(n15808), .B1(n14669), .B2(n1086), .ZN(
        n1970) );
  OAI22_X1 U2693 ( .A1(n15178), .A2(n15807), .B1(n14690), .B2(n1086), .ZN(
        n1977) );
  OAI22_X1 U2694 ( .A1(n15179), .A2(n15792), .B1(n14642), .B2(n1086), .ZN(
        n1961) );
  OAI22_X1 U2695 ( .A1(n15177), .A2(n15790), .B1(n15174), .B2(n14707), .ZN(
        n1983) );
  OAI22_X1 U2696 ( .A1(n14993), .A2(n15781), .B1(n14681), .B2(n1122), .ZN(
        n1590) );
  OAI22_X1 U2697 ( .A1(n15077), .A2(n15689), .B1(n14654), .B2(n15069), .ZN(
        n1837) );
  OAI22_X1 U2698 ( .A1(n15076), .A2(n15688), .B1(n14657), .B2(n1097), .ZN(
        n1838) );
  OAI22_X1 U2699 ( .A1(n15076), .A2(n15687), .B1(n14681), .B2(n1097), .ZN(
        n1846) );
  OAI22_X1 U2700 ( .A1(n15076), .A2(n15686), .B1(n14684), .B2(n1097), .ZN(
        n1847) );
  OAI22_X1 U2701 ( .A1(n15238), .A2(n16268), .B1(n15233), .B2(n14680), .ZN(
        n3475) );
  OAI22_X1 U2702 ( .A1(n15236), .A2(n16261), .B1(n15233), .B2(n14668), .ZN(
        n3593) );
  OAI22_X1 U2703 ( .A1(n15236), .A2(n16260), .B1(n15233), .B2(n14689), .ZN(
        n3592) );
  OAI22_X1 U2704 ( .A1(n15240), .A2(n16259), .B1(n1081), .B2(n14710), .ZN(
        n3468) );
  OAI22_X1 U2705 ( .A1(n15240), .A2(n16258), .B1(n1081), .B2(n14713), .ZN(
        n3467) );
  OAI22_X1 U2706 ( .A1(n15238), .A2(n16232), .B1(n15233), .B2(n14650), .ZN(
        n3478) );
  OAI22_X1 U2707 ( .A1(n15239), .A2(n16231), .B1(n1081), .B2(n14698), .ZN(
        n3472) );
  OAI22_X1 U2708 ( .A1(n15239), .A2(n16230), .B1(n1081), .B2(n14701), .ZN(
        n3471) );
  OAI22_X1 U2709 ( .A1(n15137), .A2(n16214), .B1(n14626), .B2(n15135), .ZN(
        n3620) );
  OAI22_X1 U2710 ( .A1(n15137), .A2(n16211), .B1(n14650), .B2(n15135), .ZN(
        n3619) );
  OAI22_X1 U2711 ( .A1(n15138), .A2(n16209), .B1(n14698), .B2(n15135), .ZN(
        n3615) );
  OAI22_X1 U2712 ( .A1(n15141), .A2(n16208), .B1(n14702), .B2(n15136), .ZN(
        n3442) );
  OAI22_X1 U2713 ( .A1(n15150), .A2(n16198), .B1(n14654), .B2(n15145), .ZN(
        n1645) );
  OAI22_X1 U2714 ( .A1(n15150), .A2(n16197), .B1(n14657), .B2(n15145), .ZN(
        n1646) );
  OAI22_X1 U2715 ( .A1(n15149), .A2(n16196), .B1(n14681), .B2(n15145), .ZN(
        n1654) );
  OAI22_X1 U2716 ( .A1(n15149), .A2(n16195), .B1(n14684), .B2(n15145), .ZN(
        n1655) );
  OAI22_X1 U2717 ( .A1(n15119), .A2(n16162), .B1(n14622), .B2(n15117), .ZN(
        n3580) );
  OAI22_X1 U2718 ( .A1(n15119), .A2(n16161), .B1(n14637), .B2(n15117), .ZN(
        n3579) );
  OAI22_X1 U2719 ( .A1(n15119), .A2(n16160), .B1(n14676), .B2(n15117), .ZN(
        n3578) );
  OAI22_X1 U2720 ( .A1(n15148), .A2(n16156), .B1(n14711), .B2(n15144), .ZN(
        n1664) );
  OAI22_X1 U2721 ( .A1(n15148), .A2(n16155), .B1(n14714), .B2(n15144), .ZN(
        n1665) );
  OAI22_X1 U2722 ( .A1(n15237), .A2(n16233), .B1(n15233), .B2(n14626), .ZN(
        n3481) );
  OAI22_X1 U2723 ( .A1(n15146), .A2(n15994), .B1(n14659), .B2(n15144), .ZN(
        n3560) );
  OAI22_X1 U2724 ( .A1(n15147), .A2(n15989), .B1(n14668), .B2(n15144), .ZN(
        n3559) );
  OAI22_X1 U2725 ( .A1(n15146), .A2(n15988), .B1(n14689), .B2(n15144), .ZN(
        n3627) );
  OAI22_X1 U2726 ( .A1(n15151), .A2(n15972), .B1(n14633), .B2(n15145), .ZN(
        n1638) );
  OAI22_X1 U2727 ( .A1(n15151), .A2(n15970), .B1(n14639), .B2(n15144), .ZN(
        n1640) );
  OAI22_X1 U2728 ( .A1(n15150), .A2(n15969), .B1(n14648), .B2(n15145), .ZN(
        n1643) );
  OAI22_X1 U2729 ( .A1(n15150), .A2(n15968), .B1(n14662), .B2(n15145), .ZN(
        n1648) );
  OAI22_X1 U2730 ( .A1(n15037), .A2(n15849), .B1(n14633), .B2(n15029), .ZN(
        n1990) );
  OAI22_X1 U2731 ( .A1(n15037), .A2(n15848), .B1(n14639), .B2(n15029), .ZN(
        n1992) );
  OAI22_X1 U2732 ( .A1(n15182), .A2(n15836), .B1(n14633), .B2(n1086), .ZN(
        n1958) );
  OAI22_X1 U2733 ( .A1(n15181), .A2(n15835), .B1(n14639), .B2(n1086), .ZN(
        n1960) );
  OAI22_X1 U2734 ( .A1(n15181), .A2(n15693), .B1(n14648), .B2(n1086), .ZN(
        n1963) );
  OAI22_X1 U2735 ( .A1(n15142), .A2(n16310), .B1(n14653), .B2(n15136), .ZN(
        n1421) );
  OAI22_X1 U2736 ( .A1(n15142), .A2(n16309), .B1(n14656), .B2(n15135), .ZN(
        n1422) );
  OAI22_X1 U2737 ( .A1(n15142), .A2(n16308), .B1(n14682), .B2(n15136), .ZN(
        n1430) );
  OAI22_X1 U2738 ( .A1(n15142), .A2(n16307), .B1(n14683), .B2(n15135), .ZN(
        n1431) );
  OAI22_X1 U2739 ( .A1(n15142), .A2(n16246), .B1(n14711), .B2(n15136), .ZN(
        n3440) );
  OAI22_X1 U2740 ( .A1(n15138), .A2(n16245), .B1(n14714), .B2(n15135), .ZN(
        n3613) );
  OAI22_X1 U2741 ( .A1(n15140), .A2(n16173), .B1(n14663), .B2(n15136), .ZN(
        n3449) );
  OAI22_X1 U2742 ( .A1(n15034), .A2(n15906), .B1(n14714), .B2(n1112), .ZN(
        n2017) );
  OAI22_X1 U2743 ( .A1(n15073), .A2(n15717), .B1(n14634), .B2(n1097), .ZN(
        n3552) );
  OAI22_X1 U2744 ( .A1(n15073), .A2(n15716), .B1(n14640), .B2(n1097), .ZN(
        n3550) );
  OAI22_X1 U2745 ( .A1(n15139), .A2(n16213), .B1(n14634), .B2(n15136), .ZN(
        n3453) );
  OAI22_X1 U2746 ( .A1(n15139), .A2(n16212), .B1(n14640), .B2(n15136), .ZN(
        n3451) );
  OAI22_X1 U2747 ( .A1(n15140), .A2(n16210), .B1(n14673), .B2(n15136), .ZN(
        n3447) );
  OAI22_X1 U2748 ( .A1(n15152), .A2(n16100), .B1(n14627), .B2(n15144), .ZN(
        n1636) );
  OAI22_X1 U2749 ( .A1(n15150), .A2(n16099), .B1(n14651), .B2(n15145), .ZN(
        n1644) );
  OAI22_X1 U2750 ( .A1(n15148), .A2(n16098), .B1(n14699), .B2(n15145), .ZN(
        n1660) );
  OAI22_X1 U2751 ( .A1(n15148), .A2(n16097), .B1(n14702), .B2(n15145), .ZN(
        n1661) );
  OAI22_X1 U2752 ( .A1(n15120), .A2(n16060), .B1(n14627), .B2(n15117), .ZN(
        n3466) );
  OAI22_X1 U2753 ( .A1(n15121), .A2(n16058), .B1(n14651), .B2(n15117), .ZN(
        n3462) );
  OAI22_X1 U2754 ( .A1(n15121), .A2(n16057), .B1(n14666), .B2(n15118), .ZN(
        n3461) );
  OAI22_X1 U2755 ( .A1(n15121), .A2(n16056), .B1(n14678), .B2(n15118), .ZN(
        n3460) );
  OAI22_X1 U2756 ( .A1(n15121), .A2(n16055), .B1(n14696), .B2(n15118), .ZN(
        n3459) );
  OAI22_X1 U2757 ( .A1(n15122), .A2(n16054), .B1(n14699), .B2(n15118), .ZN(
        n3458) );
  OAI22_X1 U2758 ( .A1(n15122), .A2(n16053), .B1(n14701), .B2(n15118), .ZN(
        n3457) );
  OAI22_X1 U2759 ( .A1(n15057), .A2(n16051), .B1(n14708), .B2(n15051), .ZN(
        n3495) );
  OAI22_X1 U2760 ( .A1(n15057), .A2(n16050), .B1(n14711), .B2(n15051), .ZN(
        n3494) );
  OAI22_X1 U2761 ( .A1(n15058), .A2(n16049), .B1(n14714), .B2(n15051), .ZN(
        n3493) );
  OAI22_X1 U2762 ( .A1(n15125), .A2(n16011), .B1(n15117), .B2(n14624), .ZN(
        n1315) );
  OAI22_X1 U2763 ( .A1(n15120), .A2(n16010), .B1(n14629), .B2(n15117), .ZN(
        n3465) );
  OAI22_X1 U2764 ( .A1(n15151), .A2(n15999), .B1(n14630), .B2(n15145), .ZN(
        n1637) );
  OAI22_X1 U2765 ( .A1(n15149), .A2(n15998), .B1(n14666), .B2(n15145), .ZN(
        n1649) );
  OAI22_X1 U2766 ( .A1(n15149), .A2(n15997), .B1(n14678), .B2(n15145), .ZN(
        n1653) );
  OAI22_X1 U2767 ( .A1(n15148), .A2(n15996), .B1(n14696), .B2(n15145), .ZN(
        n1659) );
  OAI22_X1 U2768 ( .A1(n15146), .A2(n15973), .B1(n14622), .B2(n15144), .ZN(
        n3562) );
  OAI22_X1 U2769 ( .A1(n15146), .A2(n15971), .B1(n14637), .B2(n15144), .ZN(
        n3561) );
  OAI22_X1 U2770 ( .A1(n15149), .A2(n15967), .B1(n14672), .B2(n15145), .ZN(
        n1651) );
  OAI22_X1 U2771 ( .A1(n15147), .A2(n15966), .B1(n14676), .B2(n15144), .ZN(
        n3558) );
  OAI22_X1 U2772 ( .A1(n15147), .A2(n15965), .B1(n14688), .B2(n15144), .ZN(
        n3557) );
  OAI22_X1 U2773 ( .A1(n15147), .A2(n15964), .B1(n14694), .B2(n15144), .ZN(
        n3556) );
  OAI22_X1 U2774 ( .A1(n15147), .A2(n15963), .B1(n14706), .B2(n15144), .ZN(
        n3555) );
  OAI22_X1 U2775 ( .A1(n15146), .A2(n15962), .B1(n14708), .B2(n15144), .ZN(
        n3610) );
  OAI22_X1 U2776 ( .A1(n15033), .A2(n15907), .B1(n14711), .B2(n1112), .ZN(
        n2016) );
  OAI22_X1 U2777 ( .A1(n15094), .A2(n15911), .B1(n14707), .B2(n1095), .ZN(
        n1183) );
  OAI22_X1 U2778 ( .A1(n15034), .A2(n15878), .B1(n14672), .B2(n1112), .ZN(
        n2003) );
  OAI22_X1 U2779 ( .A1(n15182), .A2(n15862), .B1(n1086), .B2(n14626), .ZN(
        n1956) );
  OAI22_X1 U2780 ( .A1(n15181), .A2(n15861), .B1(n15174), .B2(n14650), .ZN(
        n1964) );
  OAI22_X1 U2781 ( .A1(n15180), .A2(n15859), .B1(n15174), .B2(n14665), .ZN(
        n1969) );
  OAI22_X1 U2782 ( .A1(n15179), .A2(n15858), .B1(n1086), .B2(n14677), .ZN(
        n1973) );
  OAI22_X1 U2783 ( .A1(n15178), .A2(n15857), .B1(n1086), .B2(n14695), .ZN(
        n1979) );
  OAI22_X1 U2784 ( .A1(n15178), .A2(n15856), .B1(n1086), .B2(n14698), .ZN(
        n1980) );
  OAI22_X1 U2785 ( .A1(n15178), .A2(n15855), .B1(n1086), .B2(n14701), .ZN(
        n1981) );
  OAI22_X1 U2786 ( .A1(n15230), .A2(n15805), .B1(n1082), .B2(n14620), .ZN(
        n1730) );
  OAI22_X1 U2787 ( .A1(n15229), .A2(n15804), .B1(n1082), .B2(n14635), .ZN(
        n1735) );
  OAI22_X1 U2788 ( .A1(n15227), .A2(n15803), .B1(n1082), .B2(n14674), .ZN(
        n1748) );
  OAI22_X1 U2789 ( .A1(n15226), .A2(n15802), .B1(n1082), .B2(n14686), .ZN(
        n1752) );
  OAI22_X1 U2790 ( .A1(n15227), .A2(n15801), .B1(n1082), .B2(n14692), .ZN(
        n1754) );
  OAI22_X1 U2791 ( .A1(n15225), .A2(n15800), .B1(n1082), .B2(n14704), .ZN(
        n1758) );
  OAI22_X1 U2792 ( .A1(n15182), .A2(n15794), .B1(n15174), .B2(n14623), .ZN(
        n1955) );
  OAI22_X1 U2793 ( .A1(n15182), .A2(n15793), .B1(n1086), .B2(n14629), .ZN(
        n1957) );
  OAI22_X1 U2794 ( .A1(n15181), .A2(n15791), .B1(n14644), .B2(n1086), .ZN(
        n1962) );
  OAI22_X1 U2795 ( .A1(n15224), .A2(n15692), .B1(n1082), .B2(n14710), .ZN(
        n1760) );
  OAI22_X1 U2796 ( .A1(n15225), .A2(n15691), .B1(n1082), .B2(n14713), .ZN(
        n1761) );
  OAI22_X1 U2797 ( .A1(n15226), .A2(n15690), .B1(n1082), .B2(n14680), .ZN(
        n1750) );
  OAI22_X1 U2798 ( .A1(n14961), .A2(n15632), .B1(n14682), .B2(n14958), .ZN(
        n1494) );
  OAI22_X1 U2799 ( .A1(n14998), .A2(n15606), .B1(n14621), .B2(n1122), .ZN(
        n1570) );
  OAI22_X1 U2800 ( .A1(n14997), .A2(n15605), .B1(n14636), .B2(n1122), .ZN(
        n1575) );
  OAI22_X1 U2801 ( .A1(n14994), .A2(n15603), .B1(n14675), .B2(n1122), .ZN(
        n1588) );
  OAI22_X1 U2802 ( .A1(n14994), .A2(n15602), .B1(n14687), .B2(n1122), .ZN(
        n1592) );
  OAI22_X1 U2803 ( .A1(n14993), .A2(n15601), .B1(n14693), .B2(n1122), .ZN(
        n1594) );
  OAI22_X1 U2804 ( .A1(n14992), .A2(n15600), .B1(n14705), .B2(n1122), .ZN(
        n1598) );
  OAI22_X1 U2805 ( .A1(n14965), .A2(n15507), .B1(n14632), .B2(n1125), .ZN(
        n1478) );
  OAI22_X1 U2806 ( .A1(n14965), .A2(n15506), .B1(n14638), .B2(n1125), .ZN(
        n1480) );
  OAI22_X1 U2807 ( .A1(n14964), .A2(n15429), .B1(n14653), .B2(n1125), .ZN(
        n1485) );
  OAI22_X1 U2808 ( .A1(n14964), .A2(n15428), .B1(n14656), .B2(n14958), .ZN(
        n1486) );
  OAI22_X1 U2809 ( .A1(n14961), .A2(n15427), .B1(n14683), .B2(n14958), .ZN(
        n1495) );
  OAI22_X1 U2810 ( .A1(n15143), .A2(n16295), .B1(n15136), .B2(n14624), .ZN(
        n1411) );
  OAI22_X1 U2811 ( .A1(n15036), .A2(n15883), .B1(n14641), .B2(n15029), .ZN(
        n1993) );
  OAI22_X1 U2812 ( .A1(n15198), .A2(n15872), .B1(n15206), .B2(n14620), .ZN(
        n1186) );
  OAI22_X1 U2813 ( .A1(n15197), .A2(n15871), .B1(n15206), .B2(n14635), .ZN(
        n1191) );
  OAI22_X1 U2814 ( .A1(n15198), .A2(n15870), .B1(n15205), .B2(n14674), .ZN(
        n1204) );
  OAI22_X1 U2815 ( .A1(n15197), .A2(n15869), .B1(n15205), .B2(n14686), .ZN(
        n1208) );
  OAI22_X1 U2816 ( .A1(n15198), .A2(n15868), .B1(n15205), .B2(n14692), .ZN(
        n1210) );
  OAI22_X1 U2817 ( .A1(n15198), .A2(n15867), .B1(n15204), .B2(n14704), .ZN(
        n1214) );
  OAI22_X1 U2818 ( .A1(n15035), .A2(n15846), .B1(n14663), .B2(n1112), .ZN(
        n2000) );
  OAI22_X1 U2819 ( .A1(n15077), .A2(n15839), .B1(n14645), .B2(n1097), .ZN(
        n1834) );
  OAI22_X1 U2820 ( .A1(n15073), .A2(n15838), .B1(n14671), .B2(n15069), .ZN(
        n3543) );
  OAI22_X1 U2821 ( .A1(n15076), .A2(n15837), .B1(n14708), .B2(n1097), .ZN(
        n1855) );
  OAI22_X1 U2822 ( .A1(n15074), .A2(n15813), .B1(n14659), .B2(n15069), .ZN(
        n3547) );
  OAI22_X1 U2823 ( .A1(n15074), .A2(n15797), .B1(n14668), .B2(n15069), .ZN(
        n3544) );
  OAI22_X1 U2824 ( .A1(n15075), .A2(n15796), .B1(n14689), .B2(n1097), .ZN(
        n3539) );
  OAI22_X1 U2825 ( .A1(n15096), .A2(n15786), .B1(n14629), .B2(n15088), .ZN(
        n3583) );
  OAI22_X1 U2826 ( .A1(n15228), .A2(n15719), .B1(n1082), .B2(n14668), .ZN(
        n1746) );
  OAI22_X1 U2827 ( .A1(n15226), .A2(n15718), .B1(n1082), .B2(n14689), .ZN(
        n1753) );
  OAI22_X1 U2828 ( .A1(n14997), .A2(n15676), .B1(n14633), .B2(n1122), .ZN(
        n1574) );
  OAI22_X1 U2829 ( .A1(n14997), .A2(n15675), .B1(n14639), .B2(n1122), .ZN(
        n1576) );
  OAI22_X1 U2830 ( .A1(n14996), .A2(n15631), .B1(n14648), .B2(n1122), .ZN(
        n1579) );
  OAI22_X1 U2831 ( .A1(n14994), .A2(n15604), .B1(n14672), .B2(n1122), .ZN(
        n1587) );
  OAI22_X1 U2832 ( .A1(n14998), .A2(n15574), .B1(n14627), .B2(n14990), .ZN(
        n1572) );
  OAI22_X1 U2833 ( .A1(n14998), .A2(n15573), .B1(n14630), .B2(n14990), .ZN(
        n1573) );
  OAI22_X1 U2834 ( .A1(n14996), .A2(n15572), .B1(n14651), .B2(n14990), .ZN(
        n1580) );
  OAI22_X1 U2835 ( .A1(n14995), .A2(n15571), .B1(n14666), .B2(n1122), .ZN(
        n1585) );
  OAI22_X1 U2836 ( .A1(n14994), .A2(n15570), .B1(n14678), .B2(n1122), .ZN(
        n1589) );
  OAI22_X1 U2837 ( .A1(n14993), .A2(n15569), .B1(n14696), .B2(n14990), .ZN(
        n1595) );
  OAI22_X1 U2838 ( .A1(n14992), .A2(n15568), .B1(n14699), .B2(n1122), .ZN(
        n1596) );
  OAI22_X1 U2839 ( .A1(n14992), .A2(n15567), .B1(n14702), .B2(n1122), .ZN(
        n1597) );
  OAI22_X1 U2840 ( .A1(n14996), .A2(n15536), .B1(n14645), .B2(n14990), .ZN(
        n1578) );
  OAI22_X1 U2841 ( .A1(n14998), .A2(n15455), .B1(n14624), .B2(n14990), .ZN(
        n1571) );
  OAI22_X1 U2842 ( .A1(n14992), .A2(n15438), .B1(n14709), .B2(n1122), .ZN(
        n1599) );
  OAI22_X1 U2843 ( .A1(n15139), .A2(n16302), .B1(n14622), .B2(n15135), .ZN(
        n3454) );
  OAI22_X1 U2844 ( .A1(n15139), .A2(n16301), .B1(n14637), .B2(n15136), .ZN(
        n3452) );
  OAI22_X1 U2845 ( .A1(n15140), .A2(n16300), .B1(n14676), .B2(n15136), .ZN(
        n3446) );
  OAI22_X1 U2846 ( .A1(n15141), .A2(n16299), .B1(n14688), .B2(n15136), .ZN(
        n3445) );
  OAI22_X1 U2847 ( .A1(n15141), .A2(n16298), .B1(n14694), .B2(n15136), .ZN(
        n3443) );
  OAI22_X1 U2848 ( .A1(n15141), .A2(n16297), .B1(n14706), .B2(n15135), .ZN(
        n3441) );
  OAI22_X1 U2849 ( .A1(n15140), .A2(n16270), .B1(n14660), .B2(n15136), .ZN(
        n3450) );
  OAI22_X1 U2850 ( .A1(n15138), .A2(n16219), .B1(n14630), .B2(n15135), .ZN(
        n3586) );
  OAI22_X1 U2851 ( .A1(n15035), .A2(n15879), .B1(n14669), .B2(n1112), .ZN(
        n2002) );
  OAI22_X1 U2852 ( .A1(n15033), .A2(n15876), .B1(n14690), .B2(n1112), .ZN(
        n2009) );
  OAI22_X1 U2853 ( .A1(n15035), .A2(n15822), .B1(n14660), .B2(n1112), .ZN(
        n1999) );
  OAI22_X1 U2854 ( .A1(n15075), .A2(n15815), .B1(n14622), .B2(n15069), .ZN(
        n3554) );
  OAI22_X1 U2855 ( .A1(n15072), .A2(n15814), .B1(n14637), .B2(n15069), .ZN(
        n3551) );
  OAI22_X1 U2856 ( .A1(n15074), .A2(n15812), .B1(n14675), .B2(n1097), .ZN(
        n3542) );
  OAI22_X1 U2857 ( .A1(n15074), .A2(n15811), .B1(n14687), .B2(n1097), .ZN(
        n3540) );
  OAI22_X1 U2858 ( .A1(n15075), .A2(n15810), .B1(n14694), .B2(n1097), .ZN(
        n3538) );
  OAI22_X1 U2859 ( .A1(n15075), .A2(n15809), .B1(n14706), .B2(n1097), .ZN(
        n3534) );
  OAI22_X1 U2860 ( .A1(n15198), .A2(n15799), .B1(n15206), .B2(n14659), .ZN(
        n1199) );
  OAI22_X1 U2861 ( .A1(n15095), .A2(n15773), .B1(n14641), .B2(n1095), .ZN(
        n3487) );
  OAI22_X1 U2862 ( .A1(n15096), .A2(n15772), .B1(n14644), .B2(n15088), .ZN(
        n3582) );
  OAI22_X1 U2863 ( .A1(n14991), .A2(n15599), .B1(n14712), .B2(n1122), .ZN(
        n1600) );
  OAI22_X1 U2864 ( .A1(n14995), .A2(n15598), .B1(n14715), .B2(n1122), .ZN(
        n1601) );
  OAI22_X1 U2865 ( .A1(n15230), .A2(n15866), .B1(n1082), .B2(n14623), .ZN(
        n1731) );
  OAI22_X1 U2866 ( .A1(n15229), .A2(n15721), .B1(n1082), .B2(n14647), .ZN(
        n1739) );
  OAI22_X1 U2867 ( .A1(n15228), .A2(n15720), .B1(n14663), .B2(n1082), .ZN(
        n1744) );
  OAI22_X1 U2868 ( .A1(n14995), .A2(n15674), .B1(n14662), .B2(n1122), .ZN(
        n1584) );
  OAI22_X1 U2869 ( .A1(n15230), .A2(n15658), .B1(n1082), .B2(n14626), .ZN(
        n1732) );
  OAI22_X1 U2870 ( .A1(n15229), .A2(n15657), .B1(n1082), .B2(n14650), .ZN(
        n1740) );
  OAI22_X1 U2871 ( .A1(n15228), .A2(n15656), .B1(n1082), .B2(n14665), .ZN(
        n1745) );
  OAI22_X1 U2872 ( .A1(n15227), .A2(n15655), .B1(n15222), .B2(n14677), .ZN(
        n1749) );
  OAI22_X1 U2873 ( .A1(n15225), .A2(n15654), .B1(n15222), .B2(n14695), .ZN(
        n1755) );
  OAI22_X1 U2874 ( .A1(n15225), .A2(n15653), .B1(n1082), .B2(n14698), .ZN(
        n1756) );
  OAI22_X1 U2875 ( .A1(n15224), .A2(n15652), .B1(n1082), .B2(n14701), .ZN(
        n1757) );
  OAI22_X1 U2876 ( .A1(n15226), .A2(n15650), .B1(n15222), .B2(n14707), .ZN(
        n1759) );
  OAI22_X1 U2877 ( .A1(n15123), .A2(n16084), .B1(n14662), .B2(n15117), .ZN(
        n1328) );
  OAI22_X1 U2878 ( .A1(n15124), .A2(n16059), .B1(n14647), .B2(n15118), .ZN(
        n1323) );
  OAI22_X1 U2879 ( .A1(n15053), .A2(n15985), .B1(n14634), .B2(n15050), .ZN(
        n3508) );
  OAI22_X1 U2880 ( .A1(n15058), .A2(n15984), .B1(n14639), .B2(n15051), .ZN(
        n3391) );
  OAI22_X1 U2881 ( .A1(n15240), .A2(n16236), .B1(n1081), .B2(n14707), .ZN(
        n3469) );
  OAI22_X1 U2882 ( .A1(n15122), .A2(n15987), .B1(n14711), .B2(n15118), .ZN(
        n3456) );
  OAI22_X1 U2883 ( .A1(n15122), .A2(n15986), .B1(n14714), .B2(n15118), .ZN(
        n3455) );
  OAI22_X1 U2884 ( .A1(n15120), .A2(n15981), .B1(n14642), .B2(n15117), .ZN(
        n3464) );
  OAI22_X1 U2885 ( .A1(n15179), .A2(n15834), .B1(n14672), .B2(n1086), .ZN(
        n1971) );
  OAI22_X1 U2886 ( .A1(n15259), .A2(n14644), .B1(n3979), .B2(n15257), .ZN(
        n3980) );
  OAI22_X1 U2887 ( .A1(n9570), .A2(n14980), .B1(n14632), .B2(n1123), .ZN(n1542) );
  OAI22_X1 U2888 ( .A1(n9572), .A2(n14980), .B1(n14638), .B2(n1123), .ZN(n1544) );
  OAI22_X1 U2889 ( .A1(n9571), .A2(n14980), .B1(n14672), .B2(n14979), .ZN(
        n1555) );
  OAI22_X1 U2890 ( .A1(n9597), .A2(n15154), .B1(n14620), .B2(n15153), .ZN(
        n1442) );
  OAI22_X1 U2891 ( .A1(n9596), .A2(n15155), .B1(n14635), .B2(n1088), .ZN(n1447) );
  OAI22_X1 U2892 ( .A1(n3629), .A2(n15154), .B1(n14655), .B2(n1088), .ZN(n3733) );
  OAI22_X1 U2893 ( .A1(n3630), .A2(n15154), .B1(n14658), .B2(n1088), .ZN(n3732) );
  OAI22_X1 U2894 ( .A1(n9593), .A2(n15155), .B1(n14674), .B2(n1088), .ZN(n1460) );
  OAI22_X1 U2895 ( .A1(n9439), .A2(n15156), .B1(n14682), .B2(n15153), .ZN(
        n1462) );
  OAI22_X1 U2896 ( .A1(n3631), .A2(n15154), .B1(n14685), .B2(n1088), .ZN(n3731) );
  OAI22_X1 U2897 ( .A1(n9595), .A2(n15155), .B1(n14686), .B2(n1088), .ZN(n1464) );
  OAI22_X1 U2898 ( .A1(n9594), .A2(n15156), .B1(n14692), .B2(n1088), .ZN(n1466) );
  OAI22_X1 U2899 ( .A1(n9451), .A2(n15155), .B1(n14704), .B2(n1088), .ZN(n1470) );
  OAI22_X1 U2900 ( .A1(n9733), .A2(n15042), .B1(n14627), .B2(n1110), .ZN(n2020) );
  OAI22_X1 U2901 ( .A1(n9732), .A2(n15042), .B1(n14651), .B2(n1110), .ZN(n2028) );
  OAI22_X1 U2902 ( .A1(n9736), .A2(n15041), .B1(n14699), .B2(n1110), .ZN(n2044) );
  OAI22_X1 U2903 ( .A1(n9740), .A2(n15041), .B1(n14702), .B2(n15040), .ZN(
        n2045) );
  OAI22_X1 U2904 ( .A1(n9737), .A2(n15041), .B1(n14711), .B2(n1110), .ZN(n2048) );
  OAI22_X1 U2905 ( .A1(n9738), .A2(n15042), .B1(n14714), .B2(n1110), .ZN(n2049) );
  OAI22_X1 U2906 ( .A1(n9734), .A2(n15041), .B1(n14666), .B2(n1110), .ZN(n2033) );
  OAI22_X1 U2907 ( .A1(n9735), .A2(n15043), .B1(n14678), .B2(n1110), .ZN(n2037) );
  OAI22_X1 U2908 ( .A1(n9739), .A2(n15042), .B1(n14696), .B2(n15040), .ZN(
        n2043) );
  OAI22_X1 U2909 ( .A1(n3346), .A2(n15165), .B1(n14655), .B2(n15164), .ZN(
        n3744) );
  OAI22_X1 U2910 ( .A1(n3347), .A2(n15165), .B1(n14658), .B2(n1087), .ZN(n3743) );
  OAI22_X1 U2911 ( .A1(n3348), .A2(n15165), .B1(n14685), .B2(n1087), .ZN(n3739) );
  OAI22_X1 U2912 ( .A1(n9434), .A2(n15197), .B1(n15204), .B2(n14710), .ZN(
        n1216) );
  OAI22_X1 U2913 ( .A1(n9435), .A2(n15197), .B1(n15203), .B2(n14713), .ZN(
        n1217) );
  OAI22_X1 U2914 ( .A1(n3365), .A2(n15197), .B1(n14644), .B2(n15199), .ZN(
        n3754) );
  OAI22_X1 U2915 ( .A1(n3930), .A2(n15246), .B1(n15252), .B2(n14653), .ZN(
        n3937) );
  OAI22_X1 U2916 ( .A1(n3931), .A2(n15246), .B1(n15248), .B2(n14656), .ZN(
        n3936) );
  OAI22_X1 U2917 ( .A1(n3932), .A2(n15246), .B1(n15248), .B2(n14683), .ZN(
        n3935) );
  OAI22_X1 U2918 ( .A1(n3355), .A2(n15246), .B1(n15250), .B2(n14620), .ZN(
        n3764) );
  OAI22_X1 U2919 ( .A1(n3357), .A2(n15246), .B1(n15248), .B2(n14635), .ZN(
        n3763) );
  OAI22_X1 U2920 ( .A1(n3359), .A2(n15246), .B1(n15249), .B2(n14674), .ZN(
        n3761) );
  OAI22_X1 U2921 ( .A1(n3361), .A2(n15246), .B1(n15249), .B2(n14686), .ZN(
        n3759) );
  OAI22_X1 U2922 ( .A1(n3643), .A2(n15247), .B1(n15250), .B2(n14692), .ZN(
        n3758) );
  OAI22_X1 U2923 ( .A1(n3642), .A2(n15247), .B1(n15250), .B2(n14704), .ZN(
        n3757) );
  OAI22_X1 U2924 ( .A1(n3929), .A2(n15234), .B1(n1081), .B2(n14662), .ZN(n3934) );
  OAI22_X1 U2925 ( .A1(n3208), .A2(n15070), .B1(n14649), .B2(n1097), .ZN(n3549) );
  OAI22_X1 U2926 ( .A1(n3242), .A2(n15089), .B1(n14659), .B2(n1095), .ZN(n3590) );
  OAI22_X1 U2927 ( .A1(n9725), .A2(n14959), .B1(n14646), .B2(n14958), .ZN(
        n1482) );
  OAI22_X1 U2928 ( .A1(n3351), .A2(n15175), .B1(n14653), .B2(n15174), .ZN(
        n3771) );
  OAI22_X1 U2929 ( .A1(n3352), .A2(n15175), .B1(n14656), .B2(n1086), .ZN(n3770) );
  OAI22_X1 U2930 ( .A1(n9506), .A2(n15177), .B1(n14681), .B2(n1086), .ZN(n1974) );
  OAI22_X1 U2931 ( .A1(n3353), .A2(n15176), .B1(n14683), .B2(n1086), .ZN(n3768) );
  OAI22_X1 U2932 ( .A1(n9440), .A2(n15032), .B1(n14654), .B2(n1112), .ZN(n1997) );
  OAI22_X1 U2933 ( .A1(n9442), .A2(n15031), .B1(n14657), .B2(n15029), .ZN(
        n1998) );
  OAI22_X1 U2934 ( .A1(n9891), .A2(n15032), .B1(n14681), .B2(n1112), .ZN(n2006) );
  OAI22_X1 U2935 ( .A1(n9441), .A2(n15031), .B1(n14684), .B2(n1112), .ZN(n2007) );
  OAI22_X1 U2936 ( .A1(n3229), .A2(n15070), .B1(n14710), .B2(n15069), .ZN(
        n3533) );
  OAI22_X1 U2937 ( .A1(n3224), .A2(n15071), .B1(n14714), .B2(n1097), .ZN(n3532) );
  OAI22_X1 U2938 ( .A1(n3364), .A2(n15197), .B1(n15202), .B2(n14629), .ZN(
        n3755) );
  OAI22_X1 U2939 ( .A1(n7821), .A2(n15094), .B1(n14628), .B2(n1095), .ZN(n1156) );
  OAI22_X1 U2940 ( .A1(n7822), .A2(n15093), .B1(n14652), .B2(n15088), .ZN(
        n1164) );
  OAI22_X1 U2941 ( .A1(n8085), .A2(n15093), .B1(n14700), .B2(n1095), .ZN(n1180) );
  OAI22_X1 U2942 ( .A1(n8086), .A2(n15092), .B1(n14703), .B2(n1095), .ZN(n1181) );
  OAI22_X1 U2943 ( .A1(n3363), .A2(n15197), .B1(n15201), .B2(n14626), .ZN(
        n3756) );
  OAI22_X1 U2944 ( .A1(n9448), .A2(n15198), .B1(n14633), .B2(n15199), .ZN(
        n1190) );
  OAI22_X1 U2945 ( .A1(n9449), .A2(n15198), .B1(n14639), .B2(n15200), .ZN(
        n1192) );
  OAI22_X1 U2946 ( .A1(n3366), .A2(n15197), .B1(n15202), .B2(n14650), .ZN(
        n3753) );
  OAI22_X1 U2947 ( .A1(n3367), .A2(n15197), .B1(n15202), .B2(n14665), .ZN(
        n3752) );
  OAI22_X1 U2948 ( .A1(n3368), .A2(n15197), .B1(n15202), .B2(n14677), .ZN(
        n3751) );
  OAI22_X1 U2949 ( .A1(n3369), .A2(n15197), .B1(n15203), .B2(n14695), .ZN(
        n3750) );
  OAI22_X1 U2950 ( .A1(n3370), .A2(n15197), .B1(n15203), .B2(n14698), .ZN(
        n3749) );
  OAI22_X1 U2951 ( .A1(n3371), .A2(n15197), .B1(n15203), .B2(n14701), .ZN(
        n3748) );
  OAI22_X1 U2952 ( .A1(n3311), .A2(n15070), .B1(n14626), .B2(n1097), .ZN(n3553) );
  OAI22_X1 U2953 ( .A1(n3310), .A2(n15071), .B1(n14650), .B2(n1097), .ZN(n3548) );
  OAI22_X1 U2954 ( .A1(n3203), .A2(n15071), .B1(n14666), .B2(n1097), .ZN(n3545) );
  OAI22_X1 U2955 ( .A1(n3225), .A2(n15072), .B1(n14678), .B2(n1097), .ZN(n3541) );
  OAI22_X1 U2956 ( .A1(n3226), .A2(n15072), .B1(n14696), .B2(n15069), .ZN(
        n3537) );
  OAI22_X1 U2957 ( .A1(n3227), .A2(n15071), .B1(n14698), .B2(n1097), .ZN(n3536) );
  OAI22_X1 U2958 ( .A1(n3228), .A2(n15072), .B1(n14701), .B2(n1097), .ZN(n3535) );
  OAI22_X1 U2959 ( .A1(n9592), .A2(n15031), .B1(n14625), .B2(n1112), .ZN(n1987) );
  OAI22_X1 U2960 ( .A1(n9447), .A2(n15198), .B1(n14653), .B2(n15200), .ZN(
        n1197) );
  OAI22_X1 U2961 ( .A1(n9582), .A2(n15198), .B1(n14656), .B2(n15199), .ZN(
        n1198) );
  OAI22_X1 U2962 ( .A1(n9446), .A2(n15198), .B1(n14683), .B2(n15201), .ZN(
        n1207) );
  OAI22_X1 U2963 ( .A1(n3725), .A2(n15198), .B1(n15204), .B2(n14668), .ZN(
        n3780) );
  OAI22_X1 U2964 ( .A1(n3724), .A2(n15197), .B1(n15201), .B2(n14689), .ZN(
        n3779) );
  OAI22_X1 U2965 ( .A1(n3655), .A2(n15177), .B1(n1086), .B2(n14620), .ZN(n3773) );
  OAI22_X1 U2966 ( .A1(n3658), .A2(n15175), .B1(n1086), .B2(n14635), .ZN(n3772) );
  OAI22_X1 U2967 ( .A1(n3657), .A2(n15175), .B1(n1086), .B2(n14674), .ZN(n3769) );
  OAI22_X1 U2968 ( .A1(n3653), .A2(n15176), .B1(n1086), .B2(n14686), .ZN(n3767) );
  OAI22_X1 U2969 ( .A1(n3656), .A2(n15176), .B1(n1086), .B2(n14692), .ZN(n3766) );
  OAI22_X1 U2970 ( .A1(n3654), .A2(n15176), .B1(n1086), .B2(n14704), .ZN(n3765) );
  OAI22_X1 U2971 ( .A1(n3372), .A2(n15211), .B1(n15217), .B2(n14632), .ZN(
        n3785) );
  OAI22_X1 U2972 ( .A1(n3373), .A2(n15211), .B1(n15215), .B2(n14638), .ZN(
        n3784) );
  OAI22_X1 U2973 ( .A1(n3374), .A2(n15211), .B1(n15214), .B2(n14647), .ZN(
        n3783) );
  OAI22_X1 U2974 ( .A1(n3375), .A2(n15211), .B1(n14662), .B2(n15213), .ZN(
        n3782) );
  OAI22_X1 U2975 ( .A1(n3379), .A2(n15211), .B1(n15215), .B2(n14671), .ZN(
        n3781) );
  OAI22_X1 U2976 ( .A1(n3147), .A2(n15092), .B1(n14649), .B2(n1095), .ZN(n3591) );
  OAI22_X1 U2977 ( .A1(n9341), .A2(n15246), .B1(n15253), .B2(n14662), .ZN(
        n2064) );
  OAI22_X1 U2978 ( .A1(n9450), .A2(n15185), .B1(n14663), .B2(n15184), .ZN(
        n1936) );
  OAI22_X1 U2979 ( .A1(n9502), .A2(n15211), .B1(n14643), .B2(n15213), .ZN(
        n1385) );
  OAI22_X1 U2980 ( .A1(n9503), .A2(n15211), .B1(n14646), .B2(n15213), .ZN(
        n1386) );
  OAI22_X1 U2981 ( .A1(n3382), .A2(n15211), .B1(n15214), .B2(n14680), .ZN(
        n3778) );
  OAI22_X1 U2982 ( .A1(n9438), .A2(n15211), .B1(n15216), .B2(n14707), .ZN(
        n1407) );
  OAI22_X1 U2983 ( .A1(n9574), .A2(n14969), .B1(n14653), .B2(n1124), .ZN(n1517) );
  OAI22_X1 U2984 ( .A1(n9573), .A2(n14969), .B1(n14656), .B2(n14968), .ZN(
        n1518) );
  OAI22_X1 U2985 ( .A1(n9575), .A2(n14969), .B1(n14683), .B2(n1124), .ZN(n1527) );
  OAI22_X1 U2986 ( .A1(n3640), .A2(n15223), .B1(n1082), .B2(n14641), .ZN(n3786) );
  OAI22_X1 U2987 ( .A1(n3682), .A2(n15211), .B1(n15215), .B2(n14665), .ZN(
        n3737) );
  OAI22_X1 U2988 ( .A1(n3680), .A2(n15211), .B1(n15216), .B2(n14677), .ZN(
        n3736) );
  OAI22_X1 U2989 ( .A1(n3681), .A2(n15211), .B1(n15215), .B2(n14695), .ZN(
        n3735) );
  OAI22_X1 U2990 ( .A1(n9721), .A2(n15010), .B1(n14654), .B2(n1119), .ZN(n1805) );
  OAI22_X1 U2991 ( .A1(n9722), .A2(n15010), .B1(n14657), .B2(n15009), .ZN(
        n1806) );
  OAI22_X1 U2992 ( .A1(n9723), .A2(n15010), .B1(n14684), .B2(n1119), .ZN(n1815) );
  OAI22_X1 U2993 ( .A1(n9443), .A2(n15246), .B1(n15254), .B2(n14659), .ZN(
        n2063) );
  OAI22_X1 U2994 ( .A1(n9445), .A2(n15246), .B1(n15253), .B2(n14668), .ZN(
        n2066) );
  OAI22_X1 U2995 ( .A1(n9444), .A2(n15247), .B1(n15252), .B2(n14689), .ZN(
        n2073) );
  OAI22_X1 U2996 ( .A1(n3594), .A2(n15246), .B1(n15249), .B2(n14647), .ZN(
        n3762) );
  OAI22_X1 U2997 ( .A1(n3383), .A2(n15246), .B1(n15249), .B2(n14680), .ZN(
        n3760) );
  OAI22_X1 U2998 ( .A1(n9566), .A2(n15198), .B1(n14643), .B2(n15199), .ZN(
        n1193) );
  OAI22_X1 U2999 ( .A1(n9467), .A2(n14991), .B1(n14653), .B2(n1122), .ZN(n1581) );
  OAI22_X1 U3000 ( .A1(n9468), .A2(n14991), .B1(n14656), .B2(n14990), .ZN(
        n1582) );
  OAI22_X1 U3001 ( .A1(n9469), .A2(n14991), .B1(n14683), .B2(n1122), .ZN(n1591) );
  OAI22_X1 U3002 ( .A1(n9577), .A2(n15223), .B1(n15222), .B2(n14629), .ZN(
        n1733) );
  OAI22_X1 U3003 ( .A1(n9576), .A2(n15223), .B1(n14645), .B2(n15222), .ZN(
        n1738) );
  OAI22_X1 U3004 ( .A1(n8079), .A2(n15092), .B1(n14712), .B2(n15088), .ZN(
        n1184) );
  OAI22_X1 U3005 ( .A1(n8080), .A2(n15092), .B1(n14715), .B2(n1095), .ZN(n1185) );
  OAI22_X1 U3006 ( .A1(n9583), .A2(n15198), .B1(n14663), .B2(n15200), .ZN(
        n1200) );
  OAI22_X1 U3007 ( .A1(n3360), .A2(n15090), .B1(n14621), .B2(n1095), .ZN(n3491) );
  OAI22_X1 U3008 ( .A1(n3354), .A2(n15090), .B1(n14634), .B2(n1095), .ZN(n3490) );
  OAI22_X1 U3009 ( .A1(n3381), .A2(n15090), .B1(n14636), .B2(n1095), .ZN(n3489) );
  OAI22_X1 U3010 ( .A1(n3335), .A2(n15090), .B1(n14640), .B2(n1095), .ZN(n3488) );
  OAI22_X1 U3011 ( .A1(n7830), .A2(n15094), .B1(n14654), .B2(n15088), .ZN(
        n1165) );
  OAI22_X1 U3012 ( .A1(n7831), .A2(n15093), .B1(n14657), .B2(n1095), .ZN(n1166) );
  OAI22_X1 U3013 ( .A1(n3329), .A2(n15089), .B1(n14668), .B2(n1095), .ZN(n3588) );
  OAI22_X1 U3014 ( .A1(n3333), .A2(n15091), .B1(n14673), .B2(n1095), .ZN(n3486) );
  OAI22_X1 U3015 ( .A1(n3358), .A2(n15091), .B1(n14676), .B2(n1095), .ZN(n3485) );
  OAI22_X1 U3016 ( .A1(n8100), .A2(n15093), .B1(n14684), .B2(n1095), .ZN(n1175) );
  OAI22_X1 U3017 ( .A1(n3337), .A2(n15091), .B1(n14688), .B2(n1095), .ZN(n3484) );
  OAI22_X1 U3018 ( .A1(n3240), .A2(n15089), .B1(n14689), .B2(n15088), .ZN(
        n3587) );
  OAI22_X1 U3019 ( .A1(n3356), .A2(n15089), .B1(n14693), .B2(n15088), .ZN(
        n3492) );
  OAI22_X1 U3020 ( .A1(n3362), .A2(n15091), .B1(n14705), .B2(n1095), .ZN(n3483) );
  OAI22_X1 U3021 ( .A1(n9433), .A2(n15198), .B1(n14672), .B2(n15201), .ZN(
        n1203) );
  OAI22_X1 U3022 ( .A1(n9579), .A2(n15224), .B1(n14654), .B2(n15222), .ZN(
        n1741) );
  OAI22_X1 U3023 ( .A1(n9581), .A2(n15224), .B1(n14657), .B2(n15222), .ZN(
        n1742) );
  OAI22_X1 U3024 ( .A1(n9580), .A2(n15223), .B1(n14684), .B2(n1082), .ZN(n1751) );
  OAI22_X1 U3025 ( .A1(n7813), .A2(n15070), .B1(n14642), .B2(n1097), .ZN(n1833) );
  OAI22_X1 U3026 ( .A1(n9589), .A2(n15030), .B1(n14621), .B2(n1112), .ZN(n1986) );
  OAI22_X1 U3027 ( .A1(n9588), .A2(n15031), .B1(n14636), .B2(n1112), .ZN(n1991) );
  OAI22_X1 U3028 ( .A1(n9585), .A2(n15032), .B1(n14675), .B2(n1112), .ZN(n2004) );
  OAI22_X1 U3029 ( .A1(n9587), .A2(n15032), .B1(n14687), .B2(n1112), .ZN(n2008) );
  OAI22_X1 U3030 ( .A1(n9586), .A2(n15030), .B1(n14693), .B2(n1112), .ZN(n2010) );
  OAI22_X1 U3031 ( .A1(n9590), .A2(n15030), .B1(n14705), .B2(n15029), .ZN(
        n2014) );
  OAI22_X1 U3032 ( .A1(n9591), .A2(n15030), .B1(n14708), .B2(n15029), .ZN(
        n2015) );
  INV_X1 U3033 ( .A(n1107), .ZN(n15310) );
  AOI22_X1 U3034 ( .A1(n15051), .A2(n3236), .B1(Data_in[0]), .B2(n15052), .ZN(
        n1107) );
  INV_X1 U3035 ( .A(n1106), .ZN(n15309) );
  AOI22_X1 U3036 ( .A1(n15050), .A2(n3239), .B1(Data_in[5]), .B2(n15052), .ZN(
        n1106) );
  INV_X1 U3037 ( .A(n1105), .ZN(n15308) );
  AOI22_X1 U3038 ( .A1(n15051), .A2(n3243), .B1(Data_in[18]), .B2(n15052), 
        .ZN(n1105) );
  INV_X1 U3039 ( .A(n1104), .ZN(n15307) );
  AOI22_X1 U3040 ( .A1(n15050), .A2(n3244), .B1(Data_in[22]), .B2(n15052), 
        .ZN(n1104) );
  INV_X1 U3041 ( .A(n1103), .ZN(n15306) );
  AOI22_X1 U3042 ( .A1(n15051), .A2(n3258), .B1(Data_in[24]), .B2(n15053), 
        .ZN(n1103) );
  INV_X1 U3043 ( .A(n1102), .ZN(n15305) );
  AOI22_X1 U3044 ( .A1(n15050), .A2(n3245), .B1(Data_in[28]), .B2(n15053), 
        .ZN(n1102) );
  INV_X1 U3045 ( .A(Write_enable), .ZN(n16314) );
  INV_X1 U3046 ( .A(n14826), .ZN(n14812) );
endmodule


module FD_239 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_238 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_237 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_236 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_235 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_234 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_233 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_232 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_231 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_230 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_229 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_228 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_227 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_226 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_225 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_224 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_223 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_222 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_221 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_220 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_219 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_218 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_217 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_216 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_215 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_214 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_213 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_212 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_211 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_210 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_209 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_208 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_7 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_239 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_238 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_237 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_236 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_235 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_234 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_233 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_232 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_231 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_230 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_229 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_228 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_227 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_226 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_225 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_224 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_223 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_222 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_221 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_220 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_219 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_218 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_217 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_216 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_215 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_214 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_213 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_212 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_211 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_210 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_209 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_208 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FD_207 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_206 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_205 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_204 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_203 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_202 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_201 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_200 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_199 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_198 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_197 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_196 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_195 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_194 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_193 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_192 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_191 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_190 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_189 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_188 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_187 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_186 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_185 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_184 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_183 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_182 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_181 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_180 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_179 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_178 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_177 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_176 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_6 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_207 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_206 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_205 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_204 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_203 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_202 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_201 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_200 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_199 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_198 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_197 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_196 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_195 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_194 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_193 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_192 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_191 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_190 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_189 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_188 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_187 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_186 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_185 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_184 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_183 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_182 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_181 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_180 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_179 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_178 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_177 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_176 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FD_175 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_174 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_173 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_172 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_171 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_170 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_169 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_168 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_167 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_166 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_165 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_164 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_163 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_162 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_161 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_160 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_159 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_158 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_157 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_156 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_155 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_154 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_153 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_152 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_151 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_150 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_149 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_148 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_147 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_146 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_145 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_144 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_5 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_175 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_174 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_173 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_172 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_171 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_170 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_169 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_168 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_167 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_166 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_165 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_164 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_163 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_162 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_161 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_160 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_159 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_158 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_157 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_156 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_155 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_154 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_153 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_152 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_151 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_150 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_149 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_148 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_147 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_146 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_145 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_144 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FD_143 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_142 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_141 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_140 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_139 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_138 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_137 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_136 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_135 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_134 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_133 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_132 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_131 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_130 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_129 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_128 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_127 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_126 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_125 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_124 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_123 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_122 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_121 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_120 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_119 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_118 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_117 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_116 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_115 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_114 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_113 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_112 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_4 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_143 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_142 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_141 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_140 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_139 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_138 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_137 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_136 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_135 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_134 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_133 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_132 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_131 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_130 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_129 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_128 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_127 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_126 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_125 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_124 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_123 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_122 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_121 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_120 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_119 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_118 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_117 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_116 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_115 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_114 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_113 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_112 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module RDMUX ( rtype_in, itype_in, opcode_in, rd_out );
  input [4:0] rtype_in;
  input [4:0] itype_in;
  input [5:0] opcode_in;
  output [4:0] rd_out;
  wire   n7, n8, n9, n10, n11, n12, n13, n49;

  NOR4_X2 U7 ( .A1(opcode_in[2]), .A2(opcode_in[1]), .A3(opcode_in[0]), .A4(
        n13), .ZN(n8) );
  INV_X1 U2 ( .A(n8), .ZN(n49) );
  OR3_X1 U3 ( .A1(opcode_in[5]), .A2(opcode_in[4]), .A3(opcode_in[3]), .ZN(n13) );
  INV_X1 U4 ( .A(n12), .ZN(rd_out[0]) );
  AOI22_X1 U5 ( .A1(itype_in[0]), .A2(n49), .B1(rtype_in[0]), .B2(n8), .ZN(n12) );
  INV_X1 U6 ( .A(n11), .ZN(rd_out[1]) );
  AOI22_X1 U8 ( .A1(itype_in[1]), .A2(n49), .B1(rtype_in[1]), .B2(n8), .ZN(n11) );
  INV_X1 U9 ( .A(n10), .ZN(rd_out[2]) );
  AOI22_X1 U10 ( .A1(itype_in[2]), .A2(n49), .B1(rtype_in[2]), .B2(n8), .ZN(
        n10) );
  INV_X1 U11 ( .A(n9), .ZN(rd_out[3]) );
  AOI22_X1 U12 ( .A1(itype_in[3]), .A2(n49), .B1(rtype_in[3]), .B2(n8), .ZN(n9) );
  INV_X1 U13 ( .A(n7), .ZN(rd_out[4]) );
  AOI22_X1 U14 ( .A1(itype_in[4]), .A2(n49), .B1(rtype_in[4]), .B2(n8), .ZN(n7) );
endmodule


module FD_111 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_110 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_109 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_108 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_107 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT5_0 ( D, CK, RESET, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  FD_111 UFD_0 ( .D(D[0]), .CK(CK), .RESET(RESET), .Q(Q[0]) );
  FD_110 UFD_1 ( .D(D[1]), .CK(CK), .RESET(RESET), .Q(Q[1]) );
  FD_109 UFD_2 ( .D(D[2]), .CK(CK), .RESET(RESET), .Q(Q[2]) );
  FD_108 UFD_3 ( .D(D[3]), .CK(CK), .RESET(RESET), .Q(Q[3]) );
  FD_107 UFD_4 ( .D(D[4]), .CK(CK), .RESET(RESET), .Q(Q[4]) );
endmodule


module RDSELECT ( OPCODE, RD_REG_IN_RTYPE, RD_REG_IN_ITYPE, RD_OUT );
  input [5:0] OPCODE;
  input [4:0] RD_REG_IN_RTYPE;
  input [4:0] RD_REG_IN_ITYPE;
  output [4:0] RD_OUT;
  wire   n7, n8, n9, n10, n11, n12, n13, n49;

  NOR4_X2 U6 ( .A1(OPCODE[2]), .A2(OPCODE[1]), .A3(OPCODE[0]), .A4(n13), .ZN(
        n8) );
  INV_X1 U1 ( .A(n8), .ZN(n49) );
  OR3_X1 U2 ( .A1(OPCODE[5]), .A2(OPCODE[4]), .A3(OPCODE[3]), .ZN(n13) );
  INV_X1 U3 ( .A(n7), .ZN(RD_OUT[0]) );
  AOI22_X1 U4 ( .A1(RD_REG_IN_ITYPE[0]), .A2(n49), .B1(RD_REG_IN_RTYPE[0]), 
        .B2(n8), .ZN(n7) );
  INV_X1 U5 ( .A(n9), .ZN(RD_OUT[1]) );
  AOI22_X1 U7 ( .A1(RD_REG_IN_ITYPE[1]), .A2(n49), .B1(RD_REG_IN_RTYPE[1]), 
        .B2(n8), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(RD_OUT[2]) );
  AOI22_X1 U9 ( .A1(RD_REG_IN_ITYPE[2]), .A2(n49), .B1(RD_REG_IN_RTYPE[2]), 
        .B2(n8), .ZN(n10) );
  INV_X1 U10 ( .A(n11), .ZN(RD_OUT[3]) );
  AOI22_X1 U11 ( .A1(RD_REG_IN_ITYPE[3]), .A2(n49), .B1(RD_REG_IN_RTYPE[3]), 
        .B2(n8), .ZN(n11) );
  INV_X1 U12 ( .A(n12), .ZN(RD_OUT[4]) );
  AOI22_X1 U13 ( .A1(RD_REG_IN_ITYPE[4]), .A2(n49), .B1(RD_REG_IN_RTYPE[4]), 
        .B2(n8), .ZN(n12) );
endmodule


module R1_HAZARD_DETECTION ( clk, reset, OPCODE, RS1_REG_IN, RD_REG_IN, 
        TYPE_OUT, reg_one, reg_two, reg_three, alu_forwarding_one, 
        mem_forwarding_one, RS1_OUT, rs1_one, rs1_two, rs1_three );
  input [5:0] OPCODE;
  input [4:0] RS1_REG_IN;
  input [4:0] RD_REG_IN;
  output [4:0] TYPE_OUT;
  output [4:0] reg_one;
  output [4:0] reg_two;
  output [4:0] reg_three;
  output [4:0] RS1_OUT;
  output [4:0] rs1_one;
  output [4:0] rs1_two;
  output [4:0] rs1_three;
  input clk, reset;
  output alu_forwarding_one, mem_forwarding_one;
  wire   n25, n26, n31, n32, n33, n34, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n67, n68, n69,
         n70, n71, n72;

  DFFR_X1 \rd_reg_one_reg[4]  ( .D(TYPE_OUT[4]), .CK(clk), .RN(n67), .Q(
        reg_one[4]) );
  DFFR_X1 \rd_reg_one_reg[3]  ( .D(TYPE_OUT[3]), .CK(clk), .RN(n67), .Q(
        reg_one[3]) );
  DFFR_X1 \rd_reg_one_reg[2]  ( .D(TYPE_OUT[2]), .CK(clk), .RN(n67), .Q(
        reg_one[2]) );
  DFFR_X1 \rd_reg_one_reg[1]  ( .D(TYPE_OUT[1]), .CK(clk), .RN(n67), .Q(
        reg_one[1]) );
  DFFR_X1 \rd_reg_one_reg[0]  ( .D(TYPE_OUT[0]), .CK(clk), .RN(n67), .Q(
        reg_one[0]) );
  DFFR_X1 \rd_reg_two_reg[1]  ( .D(reg_one[1]), .CK(clk), .RN(n67), .Q(
        reg_two[1]), .QN(n32) );
  DFFR_X1 \rd_reg_three_reg[1]  ( .D(reg_two[1]), .CK(clk), .RN(n68), .Q(
        reg_three[1]), .QN(n34) );
  DFFR_X1 \rd_reg_two_reg[0]  ( .D(reg_one[0]), .CK(clk), .RN(n68), .Q(
        reg_two[0]), .QN(n31) );
  DFFR_X1 \rd_reg_three_reg[0]  ( .D(reg_two[0]), .CK(clk), .RN(n68), .Q(
        reg_three[0]), .QN(n33) );
  DFFR_X1 \rs1_reg_one_reg[4]  ( .D(RS1_OUT[4]), .CK(clk), .RN(n68), .Q(
        rs1_one[4]) );
  DFFR_X1 \rs1_reg_one_reg[3]  ( .D(RS1_OUT[3]), .CK(clk), .RN(n68), .Q(
        rs1_one[3]) );
  DFFR_X1 \rs1_reg_one_reg[2]  ( .D(RS1_OUT[2]), .CK(clk), .RN(n68), .Q(
        rs1_one[2]) );
  DFFR_X1 \rs1_reg_one_reg[1]  ( .D(RS1_OUT[1]), .CK(clk), .RN(n68), .Q(
        rs1_one[1]) );
  DFFR_X1 \rs1_reg_one_reg[0]  ( .D(RS1_OUT[0]), .CK(clk), .RN(n68), .Q(
        rs1_one[0]) );
  XOR2_X1 U26 ( .A(rs1_one[2]), .B(reg_three[2]), .Z(n8) );
  XOR2_X1 U27 ( .A(rs1_one[4]), .B(reg_three[4]), .Z(n7) );
  XOR2_X1 U28 ( .A(rs1_one[3]), .B(reg_three[3]), .Z(n6) );
  NAND3_X1 U29 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n5) );
  XOR2_X1 U30 ( .A(n33), .B(rs1_one[0]), .Z(n11) );
  XOR2_X1 U31 ( .A(n34), .B(rs1_one[1]), .Z(n9) );
  XOR2_X1 U32 ( .A(rs1_one[2]), .B(reg_two[2]), .Z(n15) );
  XOR2_X1 U33 ( .A(rs1_one[4]), .B(reg_two[4]), .Z(n14) );
  XOR2_X1 U34 ( .A(rs1_one[3]), .B(reg_two[3]), .Z(n13) );
  NAND3_X1 U35 ( .A1(n16), .A2(n10), .A3(n17), .ZN(n12) );
  XOR2_X1 U36 ( .A(n31), .B(rs1_one[0]), .Z(n17) );
  XOR2_X1 U37 ( .A(n32), .B(rs1_one[1]), .Z(n16) );
  OAI33_X1 U38 ( .A1(n72), .A2(OPCODE[1]), .A3(n71), .B1(n23), .B2(OPCODE[4]), 
        .B3(OPCODE[0]), .ZN(n22) );
  DFFR_X1 \rs1_reg_three_reg[4]  ( .D(rs1_two[4]), .CK(clk), .RN(n69), .Q(
        rs1_three[4]) );
  DFFR_X1 \rs1_reg_three_reg[3]  ( .D(rs1_two[3]), .CK(clk), .RN(n69), .Q(
        rs1_three[3]) );
  DFFR_X1 \rs1_reg_three_reg[2]  ( .D(rs1_two[2]), .CK(clk), .RN(n69), .Q(
        rs1_three[2]) );
  DFFR_X1 \rs1_reg_three_reg[1]  ( .D(rs1_two[1]), .CK(clk), .RN(n69), .Q(
        rs1_three[1]) );
  DFFR_X1 \rs1_reg_three_reg[0]  ( .D(rs1_two[0]), .CK(clk), .RN(n69), .Q(
        rs1_three[0]) );
  DFFR_X1 \rd_reg_two_reg[4]  ( .D(reg_one[4]), .CK(clk), .RN(n69), .Q(
        reg_two[4]) );
  DFFR_X1 \rd_reg_two_reg[3]  ( .D(reg_one[3]), .CK(clk), .RN(n69), .Q(
        reg_two[3]) );
  DFFR_X1 \rd_reg_two_reg[2]  ( .D(reg_one[2]), .CK(clk), .RN(n69), .Q(
        reg_two[2]) );
  DFFR_X1 \rd_reg_three_reg[4]  ( .D(reg_two[4]), .CK(clk), .RN(n69), .Q(
        reg_three[4]) );
  DFFR_X1 \rd_reg_three_reg[3]  ( .D(reg_two[3]), .CK(clk), .RN(n69), .Q(
        reg_three[3]) );
  DFFR_X1 \rd_reg_three_reg[2]  ( .D(reg_two[2]), .CK(clk), .RN(n69), .Q(
        reg_three[2]) );
  DFFR_X1 \rs1_reg_two_reg[2]  ( .D(rs1_one[2]), .CK(clk), .RN(n69), .Q(
        rs1_two[2]) );
  DFFR_X1 \rs1_reg_two_reg[4]  ( .D(rs1_one[4]), .CK(clk), .RN(n69), .Q(
        rs1_two[4]) );
  DFFR_X1 \rs1_reg_two_reg[3]  ( .D(rs1_one[3]), .CK(clk), .RN(n69), .Q(
        rs1_two[3]) );
  DFFR_X1 \rs1_reg_two_reg[0]  ( .D(rs1_one[0]), .CK(clk), .RN(n69), .Q(
        rs1_two[0]) );
  DFFR_X1 \rs1_reg_two_reg[1]  ( .D(rs1_one[1]), .CK(clk), .RN(n69), .Q(
        rs1_two[1]) );
  DFFR_X1 alu_forwarding_one_reg ( .D(n25), .CK(clk), .RN(n69), .Q(
        alu_forwarding_one) );
  DFFR_X1 mem_forwarding_one_reg ( .D(n26), .CK(clk), .RN(n69), .Q(
        mem_forwarding_one) );
  BUF_X1 U3 ( .A(n69), .Z(n67) );
  BUF_X1 U4 ( .A(n69), .Z(n68) );
  INV_X1 U5 ( .A(reset), .ZN(n69) );
  AND2_X1 U6 ( .A1(RD_REG_IN[0]), .A2(n19), .ZN(TYPE_OUT[0]) );
  AND2_X1 U7 ( .A1(RD_REG_IN[1]), .A2(n19), .ZN(TYPE_OUT[1]) );
  AND2_X1 U8 ( .A1(RD_REG_IN[2]), .A2(n19), .ZN(TYPE_OUT[2]) );
  AND2_X1 U9 ( .A1(RD_REG_IN[3]), .A2(n19), .ZN(TYPE_OUT[3]) );
  AND2_X1 U10 ( .A1(RD_REG_IN[4]), .A2(n19), .ZN(TYPE_OUT[4]) );
  NOR4_X1 U11 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n25) );
  NOR4_X1 U12 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n26) );
  OR4_X1 U13 ( .A1(rs1_one[3]), .A2(rs1_one[4]), .A3(rs1_one[2]), .A4(n18), 
        .ZN(n10) );
  OR2_X1 U14 ( .A1(rs1_one[1]), .A2(rs1_one[0]), .ZN(n18) );
  NOR2_X1 U15 ( .A1(OPCODE[5]), .A2(n20), .ZN(n19) );
  AOI21_X1 U16 ( .B1(OPCODE[4]), .B2(n21), .A(n22), .ZN(n20) );
  OAI21_X1 U17 ( .B1(OPCODE[2]), .B2(n72), .A(n24), .ZN(n21) );
  AND2_X1 U18 ( .A1(RS1_REG_IN[0]), .A2(n19), .ZN(RS1_OUT[0]) );
  AND2_X1 U19 ( .A1(RS1_REG_IN[1]), .A2(n19), .ZN(RS1_OUT[1]) );
  AND2_X1 U20 ( .A1(RS1_REG_IN[2]), .A2(n19), .ZN(RS1_OUT[2]) );
  AND2_X1 U21 ( .A1(RS1_REG_IN[3]), .A2(n19), .ZN(RS1_OUT[3]) );
  AND2_X1 U22 ( .A1(RS1_REG_IN[4]), .A2(n19), .ZN(RS1_OUT[4]) );
  INV_X1 U23 ( .A(OPCODE[2]), .ZN(n71) );
  INV_X1 U24 ( .A(OPCODE[3]), .ZN(n72) );
  OR3_X1 U25 ( .A1(OPCODE[0]), .A2(OPCODE[3]), .A3(n71), .ZN(n24) );
  AOI21_X1 U39 ( .B1(n70), .B2(n71), .A(OPCODE[3]), .ZN(n23) );
  INV_X1 U40 ( .A(OPCODE[1]), .ZN(n70) );
endmodule


module R2_HAZARD_DETECTION ( clk, reset, OPCODE, RS2_REG_IN, RD_REG_IN, 
        TYPE_OUT, reg_one, reg_two, reg_three, RS2_OUT, rs2_one, rs2_two, 
        rs2_three, alu_forwarding_two, mem_forwarding_two );
  input [5:0] OPCODE;
  input [4:0] RS2_REG_IN;
  input [4:0] RD_REG_IN;
  output [4:0] TYPE_OUT;
  output [4:0] reg_one;
  output [4:0] reg_two;
  output [4:0] reg_three;
  output [4:0] RS2_OUT;
  output [4:0] rs2_one;
  output [4:0] rs2_two;
  output [4:0] rs2_three;
  input clk, reset;
  output alu_forwarding_two, mem_forwarding_two;
  wire   n18, n19, n23, n24, n25, n26, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n44, n45, n46;
  assign TYPE_OUT[4] = RD_REG_IN[4];
  assign TYPE_OUT[3] = RD_REG_IN[3];
  assign TYPE_OUT[2] = RD_REG_IN[2];
  assign TYPE_OUT[1] = RD_REG_IN[1];
  assign TYPE_OUT[0] = RD_REG_IN[0];

  DFFR_X1 \rd_reg_one_reg[4]  ( .D(RD_REG_IN[4]), .CK(clk), .RN(n44), .Q(
        reg_one[4]) );
  DFFR_X1 \rd_reg_one_reg[3]  ( .D(RD_REG_IN[3]), .CK(clk), .RN(n44), .Q(
        reg_one[3]) );
  DFFR_X1 \rd_reg_one_reg[2]  ( .D(RD_REG_IN[2]), .CK(clk), .RN(n44), .Q(
        reg_one[2]) );
  DFFR_X1 \rd_reg_one_reg[1]  ( .D(RD_REG_IN[1]), .CK(clk), .RN(n44), .Q(
        reg_one[1]) );
  DFFR_X1 \rd_reg_one_reg[0]  ( .D(RD_REG_IN[0]), .CK(clk), .RN(n44), .Q(
        reg_one[0]) );
  DFFR_X1 \rd_reg_two_reg[1]  ( .D(reg_one[1]), .CK(clk), .RN(n44), .Q(
        reg_two[1]), .QN(n24) );
  DFFR_X1 \rd_reg_three_reg[1]  ( .D(reg_two[1]), .CK(clk), .RN(n45), .Q(
        reg_three[1]), .QN(n26) );
  DFFR_X1 \rd_reg_two_reg[0]  ( .D(reg_one[0]), .CK(clk), .RN(n45), .Q(
        reg_two[0]), .QN(n23) );
  DFFR_X1 \rd_reg_three_reg[0]  ( .D(reg_two[0]), .CK(clk), .RN(n45), .Q(
        reg_three[0]), .QN(n25) );
  DFFR_X1 \rs2_reg_one_reg[4]  ( .D(RS2_OUT[4]), .CK(clk), .RN(n45), .Q(
        rs2_one[4]) );
  DFFR_X1 \rs2_reg_one_reg[3]  ( .D(RS2_OUT[3]), .CK(clk), .RN(n45), .Q(
        rs2_one[3]) );
  DFFR_X1 \rs2_reg_one_reg[2]  ( .D(RS2_OUT[2]), .CK(clk), .RN(n45), .Q(
        rs2_one[2]) );
  DFFR_X1 \rs2_reg_one_reg[1]  ( .D(RS2_OUT[1]), .CK(clk), .RN(n45), .Q(
        rs2_one[1]) );
  DFFR_X1 \rs2_reg_one_reg[0]  ( .D(RS2_OUT[0]), .CK(clk), .RN(n45), .Q(
        rs2_one[0]) );
  XOR2_X1 U15 ( .A(rs2_one[2]), .B(reg_three[2]), .Z(n5) );
  XOR2_X1 U16 ( .A(rs2_one[4]), .B(reg_three[4]), .Z(n4) );
  XOR2_X1 U17 ( .A(rs2_one[3]), .B(reg_three[3]), .Z(n3) );
  NAND3_X1 U18 ( .A1(n6), .A2(n7), .A3(n8), .ZN(n2) );
  XOR2_X1 U19 ( .A(n25), .B(rs2_one[0]), .Z(n8) );
  XOR2_X1 U20 ( .A(n26), .B(rs2_one[1]), .Z(n6) );
  XOR2_X1 U21 ( .A(rs2_one[2]), .B(reg_two[2]), .Z(n12) );
  XOR2_X1 U22 ( .A(rs2_one[4]), .B(reg_two[4]), .Z(n11) );
  XOR2_X1 U23 ( .A(rs2_one[3]), .B(reg_two[3]), .Z(n10) );
  NAND3_X1 U24 ( .A1(n13), .A2(n7), .A3(n14), .ZN(n9) );
  XOR2_X1 U25 ( .A(n23), .B(rs2_one[0]), .Z(n14) );
  XOR2_X1 U26 ( .A(n24), .B(rs2_one[1]), .Z(n13) );
  DFFR_X1 \rs2_reg_three_reg[4]  ( .D(rs2_two[4]), .CK(clk), .RN(n46), .Q(
        rs2_three[4]) );
  DFFR_X1 \rs2_reg_three_reg[3]  ( .D(rs2_two[3]), .CK(clk), .RN(n46), .Q(
        rs2_three[3]) );
  DFFR_X1 \rs2_reg_three_reg[2]  ( .D(rs2_two[2]), .CK(clk), .RN(n46), .Q(
        rs2_three[2]) );
  DFFR_X1 \rs2_reg_three_reg[1]  ( .D(rs2_two[1]), .CK(clk), .RN(n46), .Q(
        rs2_three[1]) );
  DFFR_X1 \rs2_reg_three_reg[0]  ( .D(rs2_two[0]), .CK(clk), .RN(n46), .Q(
        rs2_three[0]) );
  DFFR_X1 \rd_reg_two_reg[4]  ( .D(reg_one[4]), .CK(clk), .RN(n46), .Q(
        reg_two[4]) );
  DFFR_X1 \rd_reg_two_reg[3]  ( .D(reg_one[3]), .CK(clk), .RN(n46), .Q(
        reg_two[3]) );
  DFFR_X1 \rd_reg_two_reg[2]  ( .D(reg_one[2]), .CK(clk), .RN(n46), .Q(
        reg_two[2]) );
  DFFR_X1 \rd_reg_three_reg[4]  ( .D(reg_two[4]), .CK(clk), .RN(n46), .Q(
        reg_three[4]) );
  DFFR_X1 \rd_reg_three_reg[3]  ( .D(reg_two[3]), .CK(clk), .RN(n46), .Q(
        reg_three[3]) );
  DFFR_X1 \rd_reg_three_reg[2]  ( .D(reg_two[2]), .CK(clk), .RN(n46), .Q(
        reg_three[2]) );
  DFFR_X1 \rs2_reg_two_reg[2]  ( .D(rs2_one[2]), .CK(clk), .RN(n46), .Q(
        rs2_two[2]) );
  DFFR_X1 \rs2_reg_two_reg[4]  ( .D(rs2_one[4]), .CK(clk), .RN(n46), .Q(
        rs2_two[4]) );
  DFFR_X1 \rs2_reg_two_reg[3]  ( .D(rs2_one[3]), .CK(clk), .RN(n46), .Q(
        rs2_two[3]) );
  DFFR_X1 \rs2_reg_two_reg[0]  ( .D(rs2_one[0]), .CK(clk), .RN(n46), .Q(
        rs2_two[0]) );
  DFFR_X1 \rs2_reg_two_reg[1]  ( .D(rs2_one[1]), .CK(clk), .RN(n46), .Q(
        rs2_two[1]) );
  DFFR_X1 alu_forwarding_two_reg ( .D(n18), .CK(clk), .RN(n46), .Q(
        alu_forwarding_two) );
  DFFR_X1 mem_forwarding_two_reg ( .D(n19), .CK(clk), .RN(n46), .Q(
        mem_forwarding_two) );
  BUF_X1 U3 ( .A(n46), .Z(n44) );
  BUF_X1 U4 ( .A(n46), .Z(n45) );
  INV_X1 U5 ( .A(reset), .ZN(n46) );
  NOR4_X1 U6 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n18) );
  NOR4_X1 U7 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(n19) );
  OR4_X1 U8 ( .A1(rs2_one[3]), .A2(rs2_one[4]), .A3(rs2_one[2]), .A4(n15), 
        .ZN(n7) );
  OR2_X1 U9 ( .A1(rs2_one[1]), .A2(rs2_one[0]), .ZN(n15) );
  NOR4_X1 U10 ( .A1(OPCODE[2]), .A2(OPCODE[1]), .A3(OPCODE[0]), .A4(n17), .ZN(
        n16) );
  OR3_X1 U11 ( .A1(OPCODE[5]), .A2(OPCODE[4]), .A3(OPCODE[3]), .ZN(n17) );
  AND2_X1 U12 ( .A1(RS2_REG_IN[0]), .A2(n16), .ZN(RS2_OUT[0]) );
  AND2_X1 U13 ( .A1(RS2_REG_IN[1]), .A2(n16), .ZN(RS2_OUT[1]) );
  AND2_X1 U14 ( .A1(RS2_REG_IN[2]), .A2(n16), .ZN(RS2_OUT[2]) );
  AND2_X1 U27 ( .A1(RS2_REG_IN[3]), .A2(n16), .ZN(RS2_OUT[3]) );
  AND2_X1 U28 ( .A1(RS2_REG_IN[4]), .A2(n16), .ZN(RS2_OUT[4]) );
endmodule


module HAZARD_DETECTION ( clk, reset, OPCODE, RD_REG_IN_ITYPE, RD_REG_IN_RTYPE, 
        RS1_REG_IN, RS2_REG_IN, alu_forwarding_one, mem_forwarding_one, 
        alu_forwarding_two, mem_forwarding_two, RD_OUT );
  input [5:0] OPCODE;
  input [4:0] RD_REG_IN_ITYPE;
  input [4:0] RD_REG_IN_RTYPE;
  input [4:0] RS1_REG_IN;
  input [4:0] RS2_REG_IN;
  output [4:0] RD_OUT;
  input clk, reset;
  output alu_forwarding_one, mem_forwarding_one, alu_forwarding_two,
         mem_forwarding_two;


  RDSELECT RDSEL ( .OPCODE(OPCODE), .RD_REG_IN_RTYPE(RD_REG_IN_RTYPE), 
        .RD_REG_IN_ITYPE(RD_REG_IN_ITYPE), .RD_OUT(RD_OUT) );
  R1_HAZARD_DETECTION R1_HAZARD ( .clk(clk), .reset(reset), .OPCODE(OPCODE), 
        .RS1_REG_IN(RS1_REG_IN), .RD_REG_IN(RD_OUT), .alu_forwarding_one(
        alu_forwarding_one), .mem_forwarding_one(mem_forwarding_one) );
  R2_HAZARD_DETECTION R2_HAZARD ( .clk(clk), .reset(reset), .OPCODE(OPCODE), 
        .RS2_REG_IN(RS2_REG_IN), .RD_REG_IN(RD_OUT), .alu_forwarding_two(
        alu_forwarding_two), .mem_forwarding_two(mem_forwarding_two) );
endmodule


module BOFFSET ( BOFFSET_IN, BOFFSET_OUT );
  input [15:0] BOFFSET_IN;
  output [31:0] BOFFSET_OUT;
  wire   \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[14] = BOFFSET_IN[14];
  assign BOFFSET_OUT[13] = BOFFSET_IN[13];
  assign BOFFSET_OUT[12] = BOFFSET_IN[12];
  assign BOFFSET_OUT[11] = BOFFSET_IN[11];
  assign BOFFSET_OUT[10] = BOFFSET_IN[10];
  assign BOFFSET_OUT[9] = BOFFSET_IN[9];
  assign BOFFSET_OUT[8] = BOFFSET_IN[8];
  assign BOFFSET_OUT[7] = BOFFSET_IN[7];
  assign BOFFSET_OUT[6] = BOFFSET_IN[6];
  assign BOFFSET_OUT[5] = BOFFSET_IN[5];
  assign BOFFSET_OUT[4] = BOFFSET_IN[4];
  assign BOFFSET_OUT[3] = BOFFSET_IN[3];
  assign BOFFSET_OUT[2] = BOFFSET_IN[2];
  assign BOFFSET_OUT[1] = BOFFSET_IN[1];
  assign BOFFSET_OUT[0] = BOFFSET_IN[0];
  assign BOFFSET_OUT[30] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[29] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[28] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[26] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[23] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[22] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[15] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[21] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[19] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[16] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[31] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[24] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[25] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[27] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[18] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[17] = \BOFFSET_OUT[20] ;
  assign BOFFSET_OUT[20] = \BOFFSET_OUT[20] ;

  BUF_X1 U1 ( .A(BOFFSET_IN[15]), .Z(\BOFFSET_OUT[20] ) );
endmodule


module JOFFSET ( JOFFSET_IN, JOFFSET_OUT );
  input [25:0] JOFFSET_IN;
  output [31:0] JOFFSET_OUT;

  assign JOFFSET_OUT[25] = JOFFSET_IN[25];
  assign JOFFSET_OUT[26] = JOFFSET_IN[25];
  assign JOFFSET_OUT[27] = JOFFSET_IN[25];
  assign JOFFSET_OUT[28] = JOFFSET_IN[25];
  assign JOFFSET_OUT[29] = JOFFSET_IN[25];
  assign JOFFSET_OUT[30] = JOFFSET_IN[25];
  assign JOFFSET_OUT[31] = JOFFSET_IN[25];
  assign JOFFSET_OUT[24] = JOFFSET_IN[24];
  assign JOFFSET_OUT[23] = JOFFSET_IN[23];
  assign JOFFSET_OUT[22] = JOFFSET_IN[22];
  assign JOFFSET_OUT[21] = JOFFSET_IN[21];
  assign JOFFSET_OUT[20] = JOFFSET_IN[20];
  assign JOFFSET_OUT[19] = JOFFSET_IN[19];
  assign JOFFSET_OUT[18] = JOFFSET_IN[18];
  assign JOFFSET_OUT[17] = JOFFSET_IN[17];
  assign JOFFSET_OUT[16] = JOFFSET_IN[16];
  assign JOFFSET_OUT[15] = JOFFSET_IN[15];
  assign JOFFSET_OUT[14] = JOFFSET_IN[14];
  assign JOFFSET_OUT[13] = JOFFSET_IN[13];
  assign JOFFSET_OUT[12] = JOFFSET_IN[12];
  assign JOFFSET_OUT[11] = JOFFSET_IN[11];
  assign JOFFSET_OUT[10] = JOFFSET_IN[10];
  assign JOFFSET_OUT[9] = JOFFSET_IN[9];
  assign JOFFSET_OUT[8] = JOFFSET_IN[8];
  assign JOFFSET_OUT[7] = JOFFSET_IN[7];
  assign JOFFSET_OUT[6] = JOFFSET_IN[6];
  assign JOFFSET_OUT[5] = JOFFSET_IN[5];
  assign JOFFSET_OUT[4] = JOFFSET_IN[4];
  assign JOFFSET_OUT[3] = JOFFSET_IN[3];
  assign JOFFSET_OUT[2] = JOFFSET_IN[2];
  assign JOFFSET_OUT[1] = JOFFSET_IN[1];
  assign JOFFSET_OUT[0] = JOFFSET_IN[0];

endmodule


module BRANCHDECISIONUNIT_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n33, n34, n35, n37, n38, n39,
         n40, n41, n42, n45, n46, n47, n48, n49, n50, n51, n53, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n68, n69, n70, n71, n75, n76, n77, n78,
         n79, n80, n82, n83, n85, n86, n87, n88, n89, n90, n92, n94, n96, n97,
         n98, n99, n100, n102, n104, n105, n106, n107, n108, n109, n111, n112,
         n114, n115, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n133, n134, n135, n137, n138,
         n139, n141, n142, n143, n144, n145, n146, n147, n148, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n162, n163, n165,
         n166, n167, n168, n170, n172, n173, n175, n176, n177, n178, n180,
         n181, n182, n183, n184, n185, n186, n187, n189, n190, n193, n194,
         n197, n198, n199, n201, n202, n204, n206, n207, n210, n211, n213,
         n214, n215, n217, n221, n222, n223, n226, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532;

  XOR2_X1 U197 ( .A(B[25]), .B(A[31]), .Z(n12) );
  NAND3_X1 U213 ( .A1(n82), .A2(n88), .A3(n87), .ZN(n76) );
  NAND3_X1 U221 ( .A1(n138), .A2(n137), .A3(n143), .ZN(n130) );
  OAI21_X1 U2 ( .B1(n487), .B2(n182), .A(n498), .ZN(n19) );
  OR2_X1 U3 ( .A1(n178), .A2(n226), .ZN(n193) );
  AND2_X1 U4 ( .A1(n8), .A2(n19), .ZN(n226) );
  INV_X1 U5 ( .A(n181), .ZN(n487) );
  NAND2_X1 U6 ( .A1(n498), .A2(n180), .ZN(n177) );
  NAND2_X1 U7 ( .A1(n500), .A2(n181), .ZN(n180) );
  INV_X1 U8 ( .A(n182), .ZN(n500) );
  INV_X1 U9 ( .A(n111), .ZN(n491) );
  INV_X1 U10 ( .A(n57), .ZN(n489) );
  INV_X1 U11 ( .A(n50), .ZN(n490) );
  INV_X1 U12 ( .A(n70), .ZN(n488) );
  OAI21_X1 U13 ( .B1(n222), .B2(n497), .A(n48), .ZN(n181) );
  INV_X1 U14 ( .A(n47), .ZN(n497) );
  AOI21_X1 U15 ( .B1(n65), .B2(n223), .A(n495), .ZN(n222) );
  INV_X1 U16 ( .A(n45), .ZN(n495) );
  OAI21_X1 U17 ( .B1(n482), .B2(n501), .A(n33), .ZN(n27) );
  INV_X1 U18 ( .A(n34), .ZN(n482) );
  OAI21_X1 U19 ( .B1(n483), .B2(n510), .A(n173), .ZN(n186) );
  INV_X1 U20 ( .A(n189), .ZN(n483) );
  OAI211_X1 U21 ( .C1(n519), .C2(n104), .A(n105), .B(n106), .ZN(n99) );
  INV_X1 U22 ( .A(n107), .ZN(n519) );
  AOI21_X1 U23 ( .B1(n109), .B2(n112), .A(n518), .ZN(n104) );
  NAND4_X1 U24 ( .A1(n107), .A2(n108), .A3(n109), .A4(n491), .ZN(n106) );
  OAI21_X1 U25 ( .B1(n509), .B2(n484), .A(n172), .ZN(n189) );
  INV_X1 U26 ( .A(n175), .ZN(n509) );
  INV_X1 U27 ( .A(n193), .ZN(n484) );
  OAI21_X1 U28 ( .B1(n499), .B2(n487), .A(n37), .ZN(n34) );
  INV_X1 U29 ( .A(n38), .ZN(n499) );
  OAI21_X1 U30 ( .B1(n159), .B2(n160), .A(n508), .ZN(n156) );
  NAND4_X1 U31 ( .A1(n175), .A2(n176), .A3(n167), .A4(n166), .ZN(n160) );
  INV_X1 U32 ( .A(n162), .ZN(n508) );
  AOI21_X1 U33 ( .B1(n8), .B2(n177), .A(n178), .ZN(n159) );
  OAI21_X1 U34 ( .B1(n129), .B2(n130), .A(n131), .ZN(n126) );
  NOR2_X1 U35 ( .A1(n515), .A2(n133), .ZN(n131) );
  INV_X1 U36 ( .A(n144), .ZN(n515) );
  OAI21_X1 U37 ( .B1(n527), .B2(n57), .A(n58), .ZN(n50) );
  INV_X1 U38 ( .A(n59), .ZN(n527) );
  OAI21_X1 U39 ( .B1(n75), .B2(n76), .A(n77), .ZN(n70) );
  NOR2_X1 U40 ( .A1(n11), .A2(n78), .ZN(n77) );
  AOI21_X1 U41 ( .B1(n79), .B2(n80), .A(n524), .ZN(n78) );
  AOI21_X1 U42 ( .B1(n82), .B2(n92), .A(n523), .ZN(n89) );
  INV_X1 U43 ( .A(n80), .ZN(n523) );
  AOI21_X1 U44 ( .B1(n50), .B2(n51), .A(n530), .ZN(n49) );
  INV_X1 U45 ( .A(n53), .ZN(n530) );
  OAI21_X1 U46 ( .B1(n199), .B2(n507), .A(n201), .ZN(n178) );
  INV_X1 U47 ( .A(n197), .ZN(n507) );
  AOI21_X1 U48 ( .B1(n198), .B2(n202), .A(n505), .ZN(n199) );
  INV_X1 U49 ( .A(n204), .ZN(n505) );
  NAND4_X1 U50 ( .A1(n38), .A2(n39), .A3(n26), .A4(n28), .ZN(n182) );
  AOI21_X1 U51 ( .B1(n134), .B2(n135), .A(n516), .ZN(n133) );
  INV_X1 U52 ( .A(n137), .ZN(n516) );
  NAND2_X1 U53 ( .A1(n138), .A2(n139), .ZN(n134) );
  OAI21_X1 U54 ( .B1(n513), .B2(n141), .A(n142), .ZN(n139) );
  OAI21_X1 U55 ( .B1(n485), .B2(n506), .A(n204), .ZN(n207) );
  INV_X1 U56 ( .A(n198), .ZN(n506) );
  INV_X1 U57 ( .A(n210), .ZN(n485) );
  OAI21_X1 U58 ( .B1(n163), .B2(n512), .A(n165), .ZN(n162) );
  INV_X1 U59 ( .A(n166), .ZN(n512) );
  AOI21_X1 U60 ( .B1(n167), .B2(n168), .A(n511), .ZN(n163) );
  INV_X1 U61 ( .A(n170), .ZN(n511) );
  OAI21_X1 U62 ( .B1(n504), .B2(n20), .A(n17), .ZN(n202) );
  OAI21_X1 U63 ( .B1(n501), .B2(n37), .A(n33), .ZN(n217) );
  OAI21_X1 U64 ( .B1(n510), .B2(n172), .A(n173), .ZN(n168) );
  OAI21_X1 U65 ( .B1(n494), .B2(n146), .A(n62), .ZN(n223) );
  INV_X1 U66 ( .A(n63), .ZN(n494) );
  NAND2_X1 U67 ( .A1(n111), .A2(n115), .ZN(n124) );
  NAND2_X1 U68 ( .A1(n129), .A2(n141), .ZN(n154) );
  NAND2_X1 U69 ( .A1(n75), .A2(n85), .ZN(n97) );
  NAND2_X1 U70 ( .A1(n96), .A2(n86), .ZN(n92) );
  NAND2_X1 U71 ( .A1(n87), .A2(n97), .ZN(n96) );
  NAND2_X1 U72 ( .A1(n153), .A2(n142), .ZN(n151) );
  NAND2_X1 U73 ( .A1(n143), .A2(n154), .ZN(n153) );
  NAND2_X1 U74 ( .A1(n213), .A2(n20), .ZN(n15) );
  NAND2_X1 U75 ( .A1(n19), .A2(n21), .ZN(n213) );
  NAND2_X1 U76 ( .A1(n123), .A2(n117), .ZN(n121) );
  NAND2_X1 U77 ( .A1(n108), .A2(n124), .ZN(n123) );
  NAND2_X1 U78 ( .A1(n114), .A2(n120), .ZN(n119) );
  NAND2_X1 U79 ( .A1(n109), .A2(n121), .ZN(n120) );
  NAND2_X1 U80 ( .A1(n99), .A2(n100), .ZN(n75) );
  NAND2_X1 U81 ( .A1(n126), .A2(n127), .ZN(n111) );
  NAND2_X1 U82 ( .A1(n156), .A2(n157), .ZN(n129) );
  NAND2_X1 U83 ( .A1(n24), .A2(n25), .ZN(n23) );
  NAND2_X1 U84 ( .A1(n26), .A2(n27), .ZN(n24) );
  NAND2_X1 U85 ( .A1(n185), .A2(n170), .ZN(n184) );
  NAND2_X1 U86 ( .A1(n167), .A2(n186), .ZN(n185) );
  AND2_X1 U87 ( .A1(n68), .A2(n69), .ZN(n57) );
  NAND2_X1 U88 ( .A1(n70), .A2(n71), .ZN(n68) );
  INV_X1 U89 ( .A(n176), .ZN(n510) );
  INV_X1 U90 ( .A(n39), .ZN(n501) );
  INV_X1 U91 ( .A(n16), .ZN(n504) );
  INV_X1 U92 ( .A(n214), .ZN(n498) );
  OAI21_X1 U93 ( .B1(n215), .B2(n503), .A(n29), .ZN(n214) );
  INV_X1 U94 ( .A(n28), .ZN(n503) );
  AOI21_X1 U95 ( .B1(n26), .B2(n217), .A(n502), .ZN(n215) );
  AND4_X1 U96 ( .A1(n197), .A2(n198), .A3(n16), .A4(n21), .ZN(n8) );
  INV_X1 U97 ( .A(n25), .ZN(n502) );
  INV_X1 U98 ( .A(n143), .ZN(n513) );
  OAI21_X1 U99 ( .B1(n504), .B2(n486), .A(n17), .ZN(n210) );
  INV_X1 U100 ( .A(n15), .ZN(n486) );
  OAI21_X1 U101 ( .B1(n492), .B2(n514), .A(n135), .ZN(n148) );
  INV_X1 U102 ( .A(n138), .ZN(n514) );
  INV_X1 U103 ( .A(n151), .ZN(n492) );
  OAI21_X1 U104 ( .B1(n493), .B2(n496), .A(n45), .ZN(n42) );
  INV_X1 U105 ( .A(n65), .ZN(n496) );
  INV_X1 U106 ( .A(n46), .ZN(n493) );
  OAI21_X1 U107 ( .B1(n115), .B2(n517), .A(n117), .ZN(n112) );
  INV_X1 U108 ( .A(n108), .ZN(n517) );
  NOR2_X1 U109 ( .A1(n524), .A2(n11), .ZN(n90) );
  NAND2_X1 U110 ( .A1(n61), .A2(n62), .ZN(n46) );
  NAND2_X1 U111 ( .A1(n63), .A2(n531), .ZN(n61) );
  NAND2_X1 U112 ( .A1(n114), .A2(n109), .ZN(n122) );
  INV_X1 U113 ( .A(n146), .ZN(n531) );
  NAND2_X1 U114 ( .A1(n82), .A2(n80), .ZN(n94) );
  NAND2_X1 U115 ( .A1(n65), .A2(n45), .ZN(n60) );
  NAND2_X1 U116 ( .A1(n115), .A2(n127), .ZN(n128) );
  NAND2_X1 U117 ( .A1(n86), .A2(n87), .ZN(n98) );
  NAND2_X1 U118 ( .A1(n85), .A2(n100), .ZN(n102) );
  NAND2_X1 U119 ( .A1(n135), .A2(n138), .ZN(n152) );
  NAND2_X1 U120 ( .A1(n16), .A2(n17), .ZN(n14) );
  NAND2_X1 U121 ( .A1(n39), .A2(n33), .ZN(n35) );
  NAND2_X1 U122 ( .A1(n63), .A2(n62), .ZN(n145) );
  INV_X1 U123 ( .A(n114), .ZN(n518) );
  NAND2_X1 U124 ( .A1(n26), .A2(n25), .ZN(n30) );
  NAND2_X1 U125 ( .A1(n144), .A2(n137), .ZN(n147) );
  NAND2_X1 U126 ( .A1(n141), .A2(n157), .ZN(n158) );
  NAND2_X1 U127 ( .A1(n58), .A2(n59), .ZN(n66) );
  NAND2_X1 U128 ( .A1(n204), .A2(n198), .ZN(n211) );
  NAND2_X1 U129 ( .A1(n28), .A2(n29), .ZN(n22) );
  NAND2_X1 U130 ( .A1(n142), .A2(n143), .ZN(n155) );
  INV_X1 U131 ( .A(n88), .ZN(n524) );
  NAND2_X1 U132 ( .A1(n20), .A2(n21), .ZN(n18) );
  NAND2_X1 U133 ( .A1(n37), .A2(n38), .ZN(n40) );
  NAND2_X1 U134 ( .A1(n173), .A2(n176), .ZN(n190) );
  NAND2_X1 U135 ( .A1(n201), .A2(n197), .ZN(n206) );
  NAND2_X1 U136 ( .A1(n47), .A2(n48), .ZN(n41) );
  NAND2_X1 U137 ( .A1(n170), .A2(n167), .ZN(n187) );
  NAND2_X1 U138 ( .A1(n117), .A2(n108), .ZN(n125) );
  NAND2_X1 U139 ( .A1(n172), .A2(n175), .ZN(n194) );
  NAND2_X1 U140 ( .A1(n165), .A2(n166), .ZN(n183) );
  NAND2_X1 U141 ( .A1(n105), .A2(n107), .ZN(n118) );
  AND2_X1 U142 ( .A1(n53), .A2(n51), .ZN(n9) );
  AND2_X1 U143 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U144 ( .A1(n82), .A2(n83), .ZN(n79) );
  OAI21_X1 U145 ( .B1(n520), .B2(n85), .A(n86), .ZN(n83) );
  INV_X1 U146 ( .A(n87), .ZN(n520) );
  XNOR2_X1 U147 ( .A(n89), .B(n90), .ZN(SUM[27]) );
  XNOR2_X1 U148 ( .A(n488), .B(n10), .ZN(SUM[28]) );
  XNOR2_X1 U149 ( .A(n66), .B(n489), .ZN(SUM[29]) );
  XNOR2_X1 U150 ( .A(n490), .B(n9), .ZN(SUM[30]) );
  XNOR2_X1 U151 ( .A(n49), .B(n12), .ZN(SUM[31]) );
  XNOR2_X1 U152 ( .A(n128), .B(n126), .ZN(SUM[20]) );
  XNOR2_X1 U153 ( .A(n125), .B(n124), .ZN(SUM[21]) );
  XNOR2_X1 U154 ( .A(n121), .B(n122), .ZN(SUM[22]) );
  XNOR2_X1 U155 ( .A(n99), .B(n102), .ZN(SUM[24]) );
  XNOR2_X1 U156 ( .A(n98), .B(n97), .ZN(SUM[25]) );
  XNOR2_X1 U157 ( .A(n92), .B(n94), .ZN(SUM[26]) );
  XNOR2_X1 U158 ( .A(n118), .B(n119), .ZN(SUM[23]) );
  XNOR2_X1 U159 ( .A(n211), .B(n210), .ZN(SUM[10]) );
  XNOR2_X1 U160 ( .A(n190), .B(n189), .ZN(SUM[13]) );
  XNOR2_X1 U161 ( .A(n187), .B(n186), .ZN(SUM[14]) );
  XNOR2_X1 U162 ( .A(n183), .B(n184), .ZN(SUM[15]) );
  XNOR2_X1 U163 ( .A(n158), .B(n156), .ZN(SUM[16]) );
  XNOR2_X1 U164 ( .A(n152), .B(n151), .ZN(SUM[18]) );
  XNOR2_X1 U165 ( .A(n147), .B(n148), .ZN(SUM[19]) );
  XNOR2_X1 U166 ( .A(n14), .B(n15), .ZN(SUM[9]) );
  XNOR2_X1 U167 ( .A(n155), .B(n154), .ZN(SUM[17]) );
  XNOR2_X1 U168 ( .A(n18), .B(n19), .ZN(SUM[8]) );
  XNOR2_X1 U169 ( .A(n22), .B(n23), .ZN(SUM[7]) );
  XNOR2_X1 U170 ( .A(n206), .B(n207), .ZN(SUM[11]) );
  XNOR2_X1 U171 ( .A(n194), .B(n193), .ZN(SUM[12]) );
  XNOR2_X1 U172 ( .A(n35), .B(n34), .ZN(SUM[5]) );
  XNOR2_X1 U173 ( .A(n30), .B(n27), .ZN(SUM[6]) );
  XNOR2_X1 U174 ( .A(n40), .B(n181), .ZN(SUM[4]) );
  XNOR2_X1 U175 ( .A(n60), .B(n46), .ZN(SUM[2]) );
  XNOR2_X1 U176 ( .A(n41), .B(n42), .ZN(SUM[3]) );
  AND2_X1 U177 ( .A1(n146), .A2(n221), .ZN(SUM[0]) );
  XNOR2_X1 U178 ( .A(n145), .B(n531), .ZN(SUM[1]) );
  NAND2_X1 U179 ( .A1(B[18]), .A2(A[18]), .ZN(n135) );
  NAND2_X1 U180 ( .A1(B[2]), .A2(A[2]), .ZN(n45) );
  NAND2_X1 U181 ( .A1(B[19]), .A2(A[19]), .ZN(n144) );
  NAND2_X1 U182 ( .A1(B[16]), .A2(A[16]), .ZN(n141) );
  NAND2_X1 U183 ( .A1(B[9]), .A2(A[9]), .ZN(n17) );
  NAND2_X1 U184 ( .A1(B[1]), .A2(A[1]), .ZN(n62) );
  NAND2_X1 U185 ( .A1(B[5]), .A2(A[5]), .ZN(n33) );
  NAND2_X1 U186 ( .A1(B[10]), .A2(A[10]), .ZN(n204) );
  NAND2_X1 U187 ( .A1(B[6]), .A2(A[6]), .ZN(n25) );
  NAND2_X1 U188 ( .A1(B[8]), .A2(A[8]), .ZN(n20) );
  NAND2_X1 U189 ( .A1(B[17]), .A2(A[17]), .ZN(n142) );
  NAND2_X1 U190 ( .A1(B[4]), .A2(A[4]), .ZN(n37) );
  NAND2_X1 U191 ( .A1(B[13]), .A2(A[13]), .ZN(n173) );
  NAND2_X1 U192 ( .A1(B[14]), .A2(A[14]), .ZN(n170) );
  NAND2_X1 U193 ( .A1(B[12]), .A2(A[12]), .ZN(n172) );
  OR2_X1 U194 ( .A1(B[10]), .A2(A[10]), .ZN(n198) );
  OR2_X1 U195 ( .A1(B[14]), .A2(A[14]), .ZN(n167) );
  NAND2_X1 U196 ( .A1(B[11]), .A2(A[11]), .ZN(n201) );
  OR2_X1 U198 ( .A1(B[6]), .A2(A[6]), .ZN(n26) );
  NAND2_X1 U199 ( .A1(B[0]), .A2(A[0]), .ZN(n146) );
  NAND2_X1 U200 ( .A1(B[7]), .A2(A[7]), .ZN(n29) );
  OR2_X1 U201 ( .A1(B[18]), .A2(A[18]), .ZN(n138) );
  OR2_X1 U202 ( .A1(B[17]), .A2(A[17]), .ZN(n143) );
  NAND2_X1 U203 ( .A1(B[3]), .A2(A[3]), .ZN(n48) );
  OR2_X1 U204 ( .A1(B[8]), .A2(A[8]), .ZN(n21) );
  NAND2_X1 U205 ( .A1(B[15]), .A2(A[15]), .ZN(n165) );
  OR2_X1 U206 ( .A1(B[15]), .A2(A[15]), .ZN(n166) );
  OR2_X1 U207 ( .A1(B[7]), .A2(A[7]), .ZN(n28) );
  OR2_X1 U208 ( .A1(B[11]), .A2(A[11]), .ZN(n197) );
  OR2_X1 U209 ( .A1(B[9]), .A2(A[9]), .ZN(n16) );
  OR2_X1 U210 ( .A1(B[13]), .A2(A[13]), .ZN(n176) );
  OR2_X1 U211 ( .A1(B[2]), .A2(A[2]), .ZN(n65) );
  OR2_X1 U212 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  OR2_X1 U214 ( .A1(B[4]), .A2(A[4]), .ZN(n38) );
  OR2_X1 U215 ( .A1(B[1]), .A2(A[1]), .ZN(n63) );
  OR2_X1 U216 ( .A1(B[12]), .A2(A[12]), .ZN(n175) );
  OR2_X1 U217 ( .A1(B[19]), .A2(A[19]), .ZN(n137) );
  OR2_X1 U218 ( .A1(B[16]), .A2(A[16]), .ZN(n157) );
  OR2_X1 U219 ( .A1(B[3]), .A2(A[3]), .ZN(n47) );
  NAND2_X1 U220 ( .A1(B[22]), .A2(A[22]), .ZN(n114) );
  INV_X1 U222 ( .A(B[31]), .ZN(n532) );
  NAND2_X1 U223 ( .A1(B[25]), .A2(A[30]), .ZN(n53) );
  NAND2_X1 U224 ( .A1(B[20]), .A2(A[20]), .ZN(n115) );
  NAND2_X1 U225 ( .A1(A[26]), .A2(B[29]), .ZN(n80) );
  NAND2_X1 U226 ( .A1(A[25]), .A2(B[30]), .ZN(n86) );
  NAND2_X1 U227 ( .A1(B[24]), .A2(A[24]), .ZN(n85) );
  NAND2_X1 U228 ( .A1(A[29]), .A2(B[26]), .ZN(n58) );
  NAND2_X1 U229 ( .A1(n532), .A2(n521), .ZN(n87) );
  INV_X1 U230 ( .A(A[25]), .ZN(n521) );
  NAND2_X1 U231 ( .A1(n532), .A2(n522), .ZN(n82) );
  INV_X1 U232 ( .A(A[26]), .ZN(n522) );
  OR2_X1 U233 ( .A1(B[22]), .A2(A[22]), .ZN(n109) );
  NAND2_X1 U234 ( .A1(B[21]), .A2(A[21]), .ZN(n117) );
  OR2_X1 U235 ( .A1(B[21]), .A2(A[21]), .ZN(n108) );
  NAND2_X1 U236 ( .A1(A[28]), .A2(B[27]), .ZN(n69) );
  NAND2_X1 U237 ( .A1(B[23]), .A2(A[23]), .ZN(n105) );
  NAND2_X1 U238 ( .A1(n532), .A2(n528), .ZN(n59) );
  INV_X1 U239 ( .A(A[29]), .ZN(n528) );
  OR2_X1 U240 ( .A1(B[23]), .A2(A[23]), .ZN(n107) );
  NAND2_X1 U241 ( .A1(n532), .A2(n529), .ZN(n51) );
  INV_X1 U242 ( .A(A[30]), .ZN(n529) );
  NAND2_X1 U243 ( .A1(n532), .A2(n526), .ZN(n71) );
  INV_X1 U244 ( .A(A[28]), .ZN(n526) );
  NAND2_X1 U245 ( .A1(n532), .A2(n525), .ZN(n88) );
  INV_X1 U246 ( .A(A[27]), .ZN(n525) );
  AND2_X1 U247 ( .A1(A[27]), .A2(B[28]), .ZN(n11) );
  OR2_X1 U248 ( .A1(B[20]), .A2(A[20]), .ZN(n127) );
  OR2_X1 U249 ( .A1(B[24]), .A2(A[24]), .ZN(n100) );
  OR2_X1 U250 ( .A1(B[0]), .A2(A[0]), .ZN(n221) );
endmodule


module BRANCHDECISIONUNIT_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1050, n1073, n1075, n1079, n1081, n1082, n1083, n1084, n1085, n1087,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1074, n1076, n1077, n1078, n1080, n1086, n1088, n1089, n1090,
         n1091, n1092;

  XOR2_X1 U155 ( .A(n1023), .B(n1024), .Z(SUM[9]) );
  XOR2_X1 U156 ( .A(B[7]), .B(A[7]), .Z(n1030) );
  XOR2_X1 U157 ( .A(n1031), .B(n1032), .Z(SUM[6]) );
  XOR2_X1 U158 ( .A(B[6]), .B(A[6]), .Z(n1032) );
  XOR2_X1 U159 ( .A(n1035), .B(n1036), .Z(SUM[4]) );
  XOR2_X1 U160 ( .A(B[4]), .B(A[4]), .Z(n1036) );
  XOR2_X1 U161 ( .A(n1037), .B(n1038), .Z(SUM[3]) );
  XOR2_X1 U171 ( .A(n1073), .B(n1075), .Z(SUM[21]) );
  XOR2_X1 U172 ( .A(B[26]), .B(A[21]), .Z(n1075) );
  XOR2_X1 U173 ( .A(n1081), .B(n1082), .Z(SUM[1]) );
  XOR2_X1 U174 ( .A(n1079), .B(n1084), .Z(SUM[19]) );
  XOR2_X1 U175 ( .A(B[23]), .B(A[19]), .Z(n1084) );
  XOR2_X1 U176 ( .A(n1094), .B(n1096), .Z(SUM[15]) );
  XOR2_X1 U177 ( .A(n1117), .B(n1118), .Z(SUM[11]) );
  XOR2_X1 U178 ( .A(n1119), .B(n1120), .Z(SUM[10]) );
  INV_X1 U2 ( .A(B[2]), .ZN(n1090) );
  NAND2_X1 U3 ( .A1(n1097), .A2(n1072), .ZN(n1094) );
  OAI211_X1 U4 ( .C1(n1039), .C2(n1042), .A(n1061), .B(n1040), .ZN(n1035) );
  INV_X1 U5 ( .A(n1126), .ZN(n1061) );
  AOI211_X1 U6 ( .C1(n1090), .C2(n1062), .A(n1041), .B(n1039), .ZN(n1126) );
  OAI21_X1 U7 ( .B1(n1105), .B2(n1106), .A(n1107), .ZN(n1102) );
  INV_X1 U8 ( .A(B[0]), .ZN(n1089) );
  NAND2_X1 U9 ( .A1(n1099), .A2(n1101), .ZN(n1097) );
  NOR2_X1 U10 ( .A1(n1091), .A2(n1066), .ZN(n1028) );
  OAI21_X1 U11 ( .B1(n1113), .B2(n1114), .A(n1115), .ZN(n1109) );
  AOI21_X1 U12 ( .B1(n1028), .B2(n1067), .A(n1068), .ZN(n1114) );
  INV_X1 U13 ( .A(n1025), .ZN(n1068) );
  INV_X1 U14 ( .A(B[8]), .ZN(n1091) );
  INV_X1 U15 ( .A(n1116), .ZN(n1067) );
  INV_X1 U16 ( .A(n1113), .ZN(n1070) );
  INV_X1 U17 ( .A(n1098), .ZN(n1072) );
  OAI22_X1 U18 ( .A1(n1098), .A2(n1097), .B1(n1099), .B2(n1100), .ZN(SUM[14])
         );
  AND2_X1 U19 ( .A1(n1072), .A2(n1101), .ZN(n1100) );
  NAND2_X1 U20 ( .A1(n1067), .A2(n1025), .ZN(n1023) );
  NOR2_X1 U21 ( .A1(n1069), .A2(n1113), .ZN(n1120) );
  OAI21_X1 U22 ( .B1(n1024), .B2(n1116), .A(n1025), .ZN(n1119) );
  NOR2_X1 U23 ( .A1(n1028), .A2(n1121), .ZN(n1024) );
  AOI21_X1 U24 ( .B1(n1066), .B2(n1091), .A(n1026), .ZN(n1121) );
  XNOR2_X1 U25 ( .A(n1026), .B(n1027), .ZN(SUM[8]) );
  AOI21_X1 U26 ( .B1(n1066), .B2(n1091), .A(n1028), .ZN(n1027) );
  XNOR2_X1 U27 ( .A(n1106), .B(n1108), .ZN(SUM[12]) );
  NOR2_X1 U28 ( .A1(n1105), .A2(n1071), .ZN(n1108) );
  INV_X1 U29 ( .A(n1107), .ZN(n1071) );
  XNOR2_X1 U30 ( .A(n1085), .B(n1087), .ZN(SUM[18]) );
  XNOR2_X1 U31 ( .A(B[27]), .B(n1076), .ZN(n1087) );
  NOR2_X1 U32 ( .A1(n1063), .A2(n1039), .ZN(n1038) );
  AOI22_X1 U33 ( .A1(n1041), .A2(n1042), .B1(n1062), .B2(n1090), .ZN(n1037) );
  INV_X1 U34 ( .A(n1040), .ZN(n1063) );
  XNOR2_X1 U35 ( .A(n1033), .B(n1034), .ZN(SUM[5]) );
  XNOR2_X1 U36 ( .A(B[5]), .B(n1064), .ZN(n1034) );
  INV_X1 U37 ( .A(n1115), .ZN(n1069) );
  INV_X1 U38 ( .A(A[20]), .ZN(n1077) );
  AOI211_X1 U39 ( .C1(n1109), .C2(A[11]), .A(n1065), .B(n1110), .ZN(n1106) );
  INV_X1 U40 ( .A(n1112), .ZN(n1065) );
  AOI211_X1 U41 ( .C1(n1091), .C2(n1066), .A(n1026), .B(n1111), .ZN(n1110) );
  OAI21_X1 U42 ( .B1(A[11]), .B2(n1109), .A(B[11]), .ZN(n1112) );
  OAI21_X1 U43 ( .B1(A[7]), .B2(n1058), .A(n1057), .ZN(n1026) );
  INV_X1 U44 ( .A(n1122), .ZN(n1057) );
  AOI21_X1 U45 ( .B1(n1058), .B2(A[7]), .A(B[7]), .ZN(n1122) );
  INV_X1 U46 ( .A(n1029), .ZN(n1058) );
  NOR2_X1 U47 ( .A1(A[3]), .A2(B[3]), .ZN(n1039) );
  AOI22_X1 U48 ( .A1(n1102), .A2(A[13]), .B1(n1103), .B2(B[13]), .ZN(n1099) );
  OR2_X1 U49 ( .A1(A[13]), .A2(n1102), .ZN(n1103) );
  AOI21_X1 U50 ( .B1(A[1]), .B2(B[1]), .A(n1127), .ZN(n1041) );
  NOR3_X1 U51 ( .A1(n1092), .A2(n1083), .A3(n1089), .ZN(n1127) );
  NOR2_X1 U52 ( .A1(B[1]), .A2(A[1]), .ZN(n1083) );
  AOI21_X1 U53 ( .B1(n1064), .B2(n1033), .A(n1124), .ZN(n1031) );
  AOI21_X1 U54 ( .B1(n1059), .B2(A[5]), .A(B[5]), .ZN(n1124) );
  INV_X1 U55 ( .A(n1033), .ZN(n1059) );
  NAND2_X1 U56 ( .A1(B[2]), .A2(A[2]), .ZN(n1042) );
  NAND2_X1 U57 ( .A1(B[3]), .A2(A[3]), .ZN(n1040) );
  AOI21_X1 U58 ( .B1(n1035), .B2(A[4]), .A(n1060), .ZN(n1033) );
  INV_X1 U59 ( .A(n1125), .ZN(n1060) );
  OAI21_X1 U60 ( .B1(A[4]), .B2(n1035), .A(B[4]), .ZN(n1125) );
  AOI22_X1 U61 ( .A1(n1031), .A2(A[6]), .B1(n1123), .B2(B[6]), .ZN(n1029) );
  OR2_X1 U62 ( .A1(n1031), .A2(A[6]), .ZN(n1123) );
  AND2_X1 U63 ( .A1(n1094), .A2(n1074), .ZN(n1095) );
  INV_X1 U64 ( .A(A[15]), .ZN(n1074) );
  NOR2_X1 U65 ( .A1(A[10]), .A2(B[10]), .ZN(n1113) );
  OAI211_X1 U66 ( .C1(A[11]), .C2(B[11]), .A(n1070), .B(n1067), .ZN(n1111) );
  NOR2_X1 U67 ( .A1(A[9]), .A2(B[9]), .ZN(n1116) );
  NOR2_X1 U68 ( .A1(A[14]), .A2(B[14]), .ZN(n1098) );
  NOR2_X1 U69 ( .A1(B[12]), .A2(A[12]), .ZN(n1105) );
  NAND2_X1 U70 ( .A1(B[9]), .A2(A[9]), .ZN(n1025) );
  NAND2_X1 U71 ( .A1(B[10]), .A2(A[10]), .ZN(n1115) );
  NAND2_X1 U72 ( .A1(B[12]), .A2(A[12]), .ZN(n1107) );
  NAND2_X1 U73 ( .A1(B[14]), .A2(A[14]), .ZN(n1101) );
  XNOR2_X1 U74 ( .A(B[11]), .B(A[11]), .ZN(n1118) );
  OAI21_X1 U75 ( .B1(n1069), .B2(n1119), .A(n1070), .ZN(n1117) );
  XNOR2_X1 U76 ( .A(A[15]), .B(B[15]), .ZN(n1096) );
  INV_X1 U77 ( .A(A[8]), .ZN(n1066) );
  INV_X1 U78 ( .A(A[2]), .ZN(n1062) );
  INV_X1 U79 ( .A(A[5]), .ZN(n1064) );
  XNOR2_X1 U80 ( .A(n1104), .B(n1102), .ZN(SUM[13]) );
  XNOR2_X1 U81 ( .A(A[13]), .B(B[13]), .ZN(n1104) );
  XNOR2_X1 U82 ( .A(n1029), .B(n1030), .ZN(SUM[7]) );
  INV_X1 U83 ( .A(A[0]), .ZN(n1092) );
  XNOR2_X1 U84 ( .A(n1041), .B(n1050), .ZN(SUM[2]) );
  XNOR2_X1 U85 ( .A(n1090), .B(A[2]), .ZN(n1050) );
  NOR2_X1 U86 ( .A1(n1092), .A2(n1089), .ZN(n1082) );
  AOI21_X1 U87 ( .B1(B[1]), .B2(A[1]), .A(n1083), .ZN(n1081) );
  XNOR2_X1 U88 ( .A(n1089), .B(A[0]), .ZN(SUM[0]) );
  INV_X1 U89 ( .A(A[23]), .ZN(n1078) );
  INV_X1 U90 ( .A(A[18]), .ZN(n1076) );
  INV_X1 U91 ( .A(A[25]), .ZN(n1080) );
  INV_X1 U92 ( .A(A[27]), .ZN(n1086) );
  INV_X1 U93 ( .A(A[29]), .ZN(n1088) );
  INV_X1 U94 ( .A(B[31]), .ZN(n1015) );
  OAI22_X1 U95 ( .A1(n1074), .A2(n1094), .B1(n1095), .B2(n1015), .ZN(n1016) );
  OAI222_X1 U96 ( .A1(B[31]), .A2(n1016), .B1(A[16]), .B2(B[31]), .C1(A[16]), 
        .C2(n1016), .ZN(n993) );
  INV_X1 U97 ( .A(A[17]), .ZN(n991) );
  AOI21_X1 U98 ( .B1(n991), .B2(n993), .A(n1015), .ZN(n983) );
  INV_X1 U99 ( .A(n983), .ZN(n984) );
  OAI21_X1 U100 ( .B1(n993), .B2(n991), .A(n984), .ZN(n985) );
  INV_X1 U101 ( .A(n985), .ZN(n1085) );
  OAI22_X1 U102 ( .A1(B[27]), .A2(n985), .B1(B[27]), .B2(A[18]), .ZN(n986) );
  OAI22_X1 U103 ( .A1(n1076), .A2(n986), .B1(n1085), .B2(n986), .ZN(n1079) );
  OAI21_X1 U104 ( .B1(A[19]), .B2(n1079), .A(B[23]), .ZN(n987) );
  INV_X1 U105 ( .A(n987), .ZN(n988) );
  AOI21_X1 U106 ( .B1(n1079), .B2(A[19]), .A(n988), .ZN(n995) );
  OAI21_X1 U107 ( .B1(n1077), .B2(n995), .A(n1015), .ZN(n989) );
  INV_X1 U108 ( .A(n989), .ZN(n990) );
  OAI22_X1 U109 ( .A1(n1077), .A2(n990), .B1(n995), .B2(n990), .ZN(n1073) );
  XOR2_X1 U110 ( .A(n991), .B(B[31]), .Z(n992) );
  XOR2_X1 U111 ( .A(n993), .B(n992), .Z(SUM[17]) );
  XOR2_X1 U112 ( .A(A[20]), .B(B[31]), .Z(n994) );
  XNOR2_X1 U113 ( .A(n995), .B(n994), .ZN(SUM[20]) );
  OAI21_X1 U114 ( .B1(A[21]), .B2(n1073), .A(B[26]), .ZN(n996) );
  INV_X1 U115 ( .A(n996), .ZN(n997) );
  AOI21_X1 U116 ( .B1(n1073), .B2(A[21]), .A(n997), .ZN(n1056) );
  INV_X1 U117 ( .A(n1056), .ZN(n998) );
  OAI222_X1 U118 ( .A1(B[26]), .A2(n998), .B1(A[22]), .B2(B[26]), .C1(A[22]), 
        .C2(n998), .ZN(n1019) );
  INV_X1 U119 ( .A(n1019), .ZN(n999) );
  OAI21_X1 U120 ( .B1(A[23]), .B2(n999), .A(B[23]), .ZN(n1000) );
  OAI21_X1 U121 ( .B1(n1078), .B2(n1019), .A(n1000), .ZN(n1054) );
  OR2_X1 U122 ( .A1(A[24]), .A2(n1054), .ZN(n1001) );
  AOI22_X1 U123 ( .A1(n1001), .A2(B[26]), .B1(n1054), .B2(A[24]), .ZN(n1021)
         );
  INV_X1 U124 ( .A(n1021), .ZN(n1002) );
  OAI22_X1 U125 ( .A1(B[23]), .A2(n1002), .B1(A[25]), .B2(B[23]), .ZN(n1003)
         );
  OAI22_X1 U126 ( .A1(n1080), .A2(n1003), .B1(n1021), .B2(n1003), .ZN(n1052)
         );
  OR2_X1 U127 ( .A1(A[26]), .A2(n1052), .ZN(n1004) );
  AOI22_X1 U128 ( .A1(n1004), .A2(B[26]), .B1(n1052), .B2(A[26]), .ZN(n1005)
         );
  INV_X1 U129 ( .A(n1005), .ZN(n1049) );
  OAI22_X1 U130 ( .A1(B[27]), .A2(n1049), .B1(A[27]), .B2(B[27]), .ZN(n1006)
         );
  OAI22_X1 U131 ( .A1(n1086), .A2(n1006), .B1(n1005), .B2(n1006), .ZN(n1047)
         );
  OAI21_X1 U132 ( .B1(A[28]), .B2(n1047), .A(B[23]), .ZN(n1007) );
  INV_X1 U133 ( .A(n1007), .ZN(n1008) );
  OAI22_X1 U134 ( .A1(n1008), .A2(n1047), .B1(A[28]), .B2(n1008), .ZN(n1009)
         );
  INV_X1 U135 ( .A(n1009), .ZN(n1022) );
  OAI22_X1 U136 ( .A1(B[23]), .A2(n1022), .B1(A[29]), .B2(B[23]), .ZN(n1010)
         );
  OAI22_X1 U137 ( .A1(n1088), .A2(n1010), .B1(n1010), .B2(n1009), .ZN(n1045)
         );
  OAI21_X1 U138 ( .B1(A[30]), .B2(n1045), .A(B[23]), .ZN(n1011) );
  INV_X1 U139 ( .A(n1011), .ZN(n1012) );
  OAI22_X1 U140 ( .A1(n1012), .A2(n1045), .B1(A[30]), .B2(n1012), .ZN(n1014)
         );
  XOR2_X1 U141 ( .A(n1015), .B(A[31]), .Z(n1013) );
  XOR2_X1 U142 ( .A(n1014), .B(n1013), .Z(SUM[31]) );
  XOR2_X1 U143 ( .A(A[16]), .B(n1015), .Z(n1017) );
  XNOR2_X1 U144 ( .A(n1017), .B(n1016), .ZN(SUM[16]) );
  XOR2_X1 U145 ( .A(n1078), .B(B[23]), .Z(n1018) );
  XOR2_X1 U146 ( .A(n1019), .B(n1018), .Z(SUM[23]) );
  XNOR2_X1 U147 ( .A(n1080), .B(B[23]), .ZN(n1020) );
  XNOR2_X1 U148 ( .A(n1021), .B(n1020), .ZN(SUM[25]) );
  XNOR2_X1 U149 ( .A(n1088), .B(B[23]), .ZN(n1043) );
  XOR2_X1 U150 ( .A(n1043), .B(n1022), .Z(SUM[29]) );
  XOR2_X1 U151 ( .A(A[30]), .B(B[23]), .Z(n1044) );
  XOR2_X1 U152 ( .A(n1045), .B(n1044), .Z(SUM[30]) );
  XOR2_X1 U153 ( .A(A[28]), .B(B[23]), .Z(n1046) );
  XOR2_X1 U154 ( .A(n1047), .B(n1046), .Z(SUM[28]) );
  XNOR2_X1 U162 ( .A(n1086), .B(B[27]), .ZN(n1048) );
  XOR2_X1 U163 ( .A(n1049), .B(n1048), .Z(SUM[27]) );
  XOR2_X1 U164 ( .A(A[26]), .B(B[26]), .Z(n1051) );
  XOR2_X1 U165 ( .A(n1052), .B(n1051), .Z(SUM[26]) );
  XOR2_X1 U166 ( .A(A[24]), .B(B[26]), .Z(n1053) );
  XOR2_X1 U167 ( .A(n1054), .B(n1053), .Z(SUM[24]) );
  XOR2_X1 U168 ( .A(A[22]), .B(B[26]), .Z(n1055) );
  XNOR2_X1 U169 ( .A(n1056), .B(n1055), .ZN(SUM[22]) );
endmodule


module BRANCHDECISIONUNIT_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1003, n1004, n1005, n1006, n1013, n1014, n1063, n1067, n1069,
         n1075, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n1002, n1007, n1008, n1009,
         n1010, n1011, n1012, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1064, n1065, n1066, n1068, n1070, n1071, n1072, n1073, n1074,
         n1076, n1077, n1117, n1118, n1120, n1121;

  XOR2_X1 U179 ( .A(n981), .B(n982), .Z(SUM[9]) );
  XOR2_X1 U180 ( .A(n984), .B(n985), .Z(SUM[8]) );
  XOR2_X1 U181 ( .A(n987), .B(n988), .Z(SUM[7]) );
  XOR2_X1 U182 ( .A(B[7]), .B(A[7]), .Z(n988) );
  XOR2_X1 U183 ( .A(n992), .B(n990), .Z(SUM[6]) );
  XOR2_X1 U184 ( .A(n999), .B(n1000), .Z(SUM[5]) );
  XOR2_X1 U205 ( .A(n1118), .B(n1063), .Z(SUM[1]) );
  XOR2_X1 U206 ( .A(B[1]), .B(A[1]), .Z(n1063) );
  XOR2_X1 U209 ( .A(n1069), .B(n1067), .Z(SUM[18]) );
  XOR2_X1 U211 ( .A(n1085), .B(n1086), .Z(SUM[15]) );
  XOR2_X1 U212 ( .A(n1073), .B(B[17]), .Z(n1085) );
  XOR2_X1 U213 ( .A(n1087), .B(n1089), .Z(SUM[14]) );
  XOR2_X1 U214 ( .A(n1090), .B(n1091), .Z(SUM[13]) );
  XOR2_X1 U215 ( .A(n1083), .B(n1093), .Z(SUM[12]) );
  NAND3_X1 U216 ( .A1(n984), .A2(n1062), .A3(n1096), .ZN(n1095) );
  XOR2_X1 U217 ( .A(n1103), .B(n1104), .Z(SUM[11]) );
  XOR2_X1 U218 ( .A(n1121), .B(A[11]), .Z(n1103) );
  INV_X1 U2 ( .A(n941), .ZN(n940) );
  INV_X1 U3 ( .A(B[31]), .ZN(n941) );
  OAI221_X1 U4 ( .B1(n1110), .B2(n1120), .C1(n991), .C2(n1061), .A(n1111), 
        .ZN(n984) );
  INV_X1 U5 ( .A(B[7]), .ZN(n1120) );
  AND2_X1 U6 ( .A1(n991), .A2(n1061), .ZN(n1110) );
  OAI211_X1 U7 ( .C1(n1001), .C2(n1112), .A(n1060), .B(n1059), .ZN(n1111) );
  NOR2_X1 U8 ( .A1(n1054), .A2(n998), .ZN(n1001) );
  AOI21_X1 U9 ( .B1(n1068), .B2(n1083), .A(n1084), .ZN(n1080) );
  AOI21_X1 U10 ( .B1(n1066), .B2(n1121), .A(n1097), .ZN(n1096) );
  INV_X1 U11 ( .A(B[11]), .ZN(n1121) );
  INV_X1 U12 ( .A(n989), .ZN(n1060) );
  INV_X1 U13 ( .A(n1092), .ZN(n1068) );
  INV_X1 U14 ( .A(n980), .ZN(n1118) );
  NAND2_X1 U15 ( .A1(n1003), .A2(n993), .ZN(n1112) );
  INV_X1 U16 ( .A(n1098), .ZN(n1064) );
  INV_X1 U17 ( .A(n1088), .ZN(n1071) );
  INV_X1 U18 ( .A(n986), .ZN(n1062) );
  INV_X1 U19 ( .A(n1114), .ZN(n1054) );
  OAI21_X1 U20 ( .B1(n997), .B2(n1004), .A(n1006), .ZN(n1114) );
  NAND2_X1 U21 ( .A1(n991), .A2(n1060), .ZN(n992) );
  XNOR2_X1 U22 ( .A(n939), .B(n1054), .ZN(SUM[4]) );
  NOR2_X1 U23 ( .A1(n998), .A2(n1058), .ZN(n939) );
  NAND2_X1 U24 ( .A1(n1070), .A2(n1081), .ZN(n1091) );
  INV_X1 U25 ( .A(n1079), .ZN(n1070) );
  NOR2_X1 U26 ( .A1(n1088), .A2(n1072), .ZN(n1089) );
  NOR2_X1 U27 ( .A1(n1084), .A2(n1092), .ZN(n1093) );
  AOI21_X1 U28 ( .B1(n1087), .B2(n1071), .A(n1072), .ZN(n1086) );
  OAI21_X1 U29 ( .B1(n1079), .B2(n1090), .A(n1081), .ZN(n1087) );
  OAI21_X1 U30 ( .B1(n1084), .B2(n1083), .A(n1068), .ZN(n1090) );
  AOI21_X1 U31 ( .B1(n981), .B2(n983), .A(n1097), .ZN(n1105) );
  XNOR2_X1 U32 ( .A(n1004), .B(n1005), .ZN(SUM[3]) );
  NOR2_X1 U33 ( .A1(n1057), .A2(n997), .ZN(n1005) );
  XNOR2_X1 U34 ( .A(n1053), .B(n1075), .ZN(SUM[16]) );
  INV_X1 U35 ( .A(n1003), .ZN(n1058) );
  INV_X1 U36 ( .A(n1082), .ZN(n1072) );
  INV_X1 U37 ( .A(n1006), .ZN(n1057) );
  OAI22_X1 U38 ( .A1(B[9]), .A2(A[9]), .B1(B[10]), .B2(A[10]), .ZN(n1097) );
  OAI221_X1 U39 ( .B1(n1097), .B2(n1100), .C1(n1101), .C2(n983), .A(n1102), 
        .ZN(n1098) );
  NOR2_X1 U40 ( .A1(A[10]), .A2(B[10]), .ZN(n1101) );
  NAND2_X1 U41 ( .A1(B[8]), .A2(A[8]), .ZN(n1100) );
  NOR2_X1 U42 ( .A1(A[3]), .A2(B[3]), .ZN(n997) );
  NOR2_X1 U43 ( .A1(A[13]), .A2(B[13]), .ZN(n1079) );
  AOI21_X1 U44 ( .B1(A[2]), .B2(B[2]), .A(n1055), .ZN(n1004) );
  NOR2_X1 U45 ( .A1(A[4]), .A2(B[4]), .ZN(n998) );
  OAI21_X1 U46 ( .B1(n980), .B2(n1056), .A(n1116), .ZN(n1014) );
  INV_X1 U47 ( .A(A[1]), .ZN(n1056) );
  OAI21_X1 U48 ( .B1(n1118), .B2(A[1]), .A(B[1]), .ZN(n1116) );
  INV_X1 U49 ( .A(A[30]), .ZN(n1117) );
  NOR2_X1 U50 ( .A1(A[14]), .A2(B[14]), .ZN(n1088) );
  NOR2_X1 U51 ( .A1(A[8]), .A2(B[8]), .ZN(n986) );
  NOR2_X1 U52 ( .A1(A[6]), .A2(B[6]), .ZN(n989) );
  INV_X1 U53 ( .A(n1115), .ZN(n1055) );
  OAI21_X1 U54 ( .B1(B[2]), .B2(A[2]), .A(n1014), .ZN(n1115) );
  NOR2_X1 U55 ( .A1(B[12]), .A2(A[12]), .ZN(n1092) );
  NAND2_X1 U56 ( .A1(B[9]), .A2(A[9]), .ZN(n983) );
  INV_X1 U57 ( .A(A[28]), .ZN(n1077) );
  INV_X1 U58 ( .A(A[23]), .ZN(n1074) );
  NAND2_X1 U59 ( .A1(B[6]), .A2(A[6]), .ZN(n991) );
  NAND2_X1 U60 ( .A1(B[10]), .A2(A[10]), .ZN(n1102) );
  NAND2_X1 U61 ( .A1(B[13]), .A2(A[13]), .ZN(n1081) );
  NAND2_X1 U62 ( .A1(B[5]), .A2(A[5]), .ZN(n993) );
  NAND2_X1 U63 ( .A1(B[0]), .A2(A[0]), .ZN(n980) );
  NAND2_X1 U64 ( .A1(n1094), .A2(n1095), .ZN(n1083) );
  OAI21_X1 U65 ( .B1(A[11]), .B2(n1098), .A(n1099), .ZN(n1094) );
  OAI21_X1 U66 ( .B1(n1064), .B2(n1066), .A(n1121), .ZN(n1099) );
  NAND2_X1 U67 ( .A1(B[4]), .A2(A[4]), .ZN(n1003) );
  NAND2_X1 U68 ( .A1(B[14]), .A2(A[14]), .ZN(n1082) );
  NAND2_X1 U69 ( .A1(B[3]), .A2(A[3]), .ZN(n1006) );
  OAI211_X1 U70 ( .C1(n1079), .C2(n1080), .A(n1081), .B(n1082), .ZN(n1078) );
  AND2_X1 U71 ( .A1(B[12]), .A2(A[12]), .ZN(n1084) );
  INV_X1 U72 ( .A(n1113), .ZN(n1059) );
  OAI22_X1 U73 ( .A1(A[5]), .A2(B[5]), .B1(A[7]), .B2(B[7]), .ZN(n1113) );
  OAI21_X1 U74 ( .B1(n1109), .B2(n984), .A(n1062), .ZN(n981) );
  AND2_X1 U75 ( .A1(A[8]), .A2(B[8]), .ZN(n1109) );
  OAI21_X1 U76 ( .B1(B[9]), .B2(A[9]), .A(n983), .ZN(n982) );
  OAI21_X1 U77 ( .B1(n989), .B2(n990), .A(n991), .ZN(n987) );
  OAI21_X1 U78 ( .B1(B[5]), .B2(A[5]), .A(n993), .ZN(n999) );
  NOR2_X1 U79 ( .A1(n1001), .A2(n1058), .ZN(n1000) );
  NOR2_X1 U80 ( .A1(n1105), .A2(n1065), .ZN(n1104) );
  INV_X1 U81 ( .A(n1102), .ZN(n1065) );
  AOI21_X1 U82 ( .B1(B[8]), .B2(A[8]), .A(n986), .ZN(n985) );
  XNOR2_X1 U83 ( .A(n1013), .B(n1014), .ZN(SUM[2]) );
  XNOR2_X1 U84 ( .A(A[2]), .B(B[2]), .ZN(n1013) );
  XNOR2_X1 U85 ( .A(n1106), .B(n1107), .ZN(SUM[10]) );
  OAI21_X1 U86 ( .B1(A[10]), .B2(B[10]), .A(n1102), .ZN(n1107) );
  OAI21_X1 U87 ( .B1(n1108), .B2(n981), .A(n983), .ZN(n1106) );
  NOR2_X1 U88 ( .A1(A[9]), .A2(B[9]), .ZN(n1108) );
  AND2_X1 U89 ( .A1(n993), .A2(n994), .ZN(n990) );
  OAI22_X1 U90 ( .A1(A[5]), .A2(B[5]), .B1(n995), .B2(n1058), .ZN(n994) );
  NOR3_X1 U91 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
  AOI211_X1 U92 ( .C1(B[2]), .C2(A[2]), .A(n1057), .B(n1055), .ZN(n996) );
  INV_X1 U93 ( .A(A[11]), .ZN(n1066) );
  INV_X1 U94 ( .A(n979), .ZN(SUM[0]) );
  OAI21_X1 U95 ( .B1(B[0]), .B2(A[0]), .A(n980), .ZN(n979) );
  INV_X1 U96 ( .A(A[7]), .ZN(n1061) );
  INV_X1 U97 ( .A(A[15]), .ZN(n1073) );
  INV_X1 U98 ( .A(A[24]), .ZN(n1076) );
  NOR2_X1 U99 ( .A1(B[22]), .A2(A[20]), .ZN(n1033) );
  NOR2_X1 U100 ( .A1(n940), .A2(A[18]), .ZN(n1038) );
  INV_X1 U101 ( .A(B[17]), .ZN(n1041) );
  OAI211_X1 U102 ( .C1(A[15]), .C2(B[17]), .A(n1078), .B(n1071), .ZN(n942) );
  OAI21_X1 U103 ( .B1(n1073), .B2(n1041), .A(n942), .ZN(n943) );
  INV_X1 U104 ( .A(n943), .ZN(n1053) );
  NOR2_X1 U105 ( .A1(A[16]), .A2(B[22]), .ZN(n1048) );
  NAND2_X1 U106 ( .A1(A[16]), .A2(B[22]), .ZN(n1046) );
  OAI21_X1 U107 ( .B1(n1053), .B2(n1048), .A(n1046), .ZN(n1042) );
  OAI21_X1 U108 ( .B1(A[17]), .B2(n1042), .A(B[17]), .ZN(n944) );
  INV_X1 U109 ( .A(n944), .ZN(n945) );
  OAI22_X1 U110 ( .A1(n945), .A2(n1042), .B1(A[17]), .B2(n945), .ZN(n1067) );
  NOR2_X1 U111 ( .A1(n1038), .A2(n1067), .ZN(n946) );
  NOR2_X1 U112 ( .A1(n940), .A2(n946), .ZN(n948) );
  INV_X1 U113 ( .A(A[19]), .ZN(n947) );
  INV_X1 U114 ( .A(n946), .ZN(n1009) );
  NAND2_X1 U115 ( .A1(A[18]), .A2(n940), .ZN(n1040) );
  OAI221_X1 U116 ( .B1(n948), .B2(n947), .C1(n941), .C2(n1009), .A(n1040), 
        .ZN(n951) );
  NAND2_X1 U117 ( .A1(A[20]), .A2(B[22]), .ZN(n963) );
  INV_X1 U118 ( .A(n963), .ZN(n960) );
  NOR2_X1 U119 ( .A1(n951), .A2(n960), .ZN(n1034) );
  INV_X1 U120 ( .A(n1034), .ZN(n950) );
  OAI21_X1 U121 ( .B1(n1033), .B2(n960), .A(n951), .ZN(n949) );
  OAI21_X1 U122 ( .B1(n1033), .B2(n950), .A(n949), .ZN(SUM[20]) );
  INV_X1 U123 ( .A(A[21]), .ZN(n1035) );
  AOI21_X1 U124 ( .B1(n1035), .B2(n941), .A(n1033), .ZN(n952) );
  NAND2_X1 U125 ( .A1(n952), .A2(n951), .ZN(n962) );
  NAND2_X1 U126 ( .A1(A[22]), .A2(B[22]), .ZN(n959) );
  NAND2_X1 U127 ( .A1(n962), .A2(n959), .ZN(n955) );
  INV_X1 U128 ( .A(n952), .ZN(n953) );
  OAI22_X1 U129 ( .A1(n1035), .A2(n941), .B1(n953), .B2(n963), .ZN(n954) );
  NOR2_X1 U130 ( .A1(A[22]), .A2(B[22]), .ZN(n1049) );
  INV_X1 U131 ( .A(n1049), .ZN(n964) );
  OAI21_X1 U132 ( .B1(n955), .B2(n954), .A(n964), .ZN(n956) );
  XOR2_X1 U133 ( .A(n941), .B(n956), .Z(n958) );
  XOR2_X1 U134 ( .A(n956), .B(n940), .Z(n957) );
  OAI22_X1 U135 ( .A1(n1074), .A2(n958), .B1(A[23]), .B2(n957), .ZN(SUM[23])
         );
  NOR2_X1 U136 ( .A1(n940), .A2(A[26]), .ZN(n975) );
  NOR2_X1 U137 ( .A1(n940), .A2(A[25]), .ZN(n1015) );
  NOR3_X1 U138 ( .A1(n975), .A2(n1076), .A3(n1015), .ZN(n968) );
  INV_X1 U139 ( .A(n959), .ZN(n1050) );
  OAI21_X1 U140 ( .B1(B[30]), .B2(n960), .A(A[21]), .ZN(n961) );
  OAI211_X1 U141 ( .C1(n941), .C2(n963), .A(n962), .B(n961), .ZN(n1052) );
  OAI21_X1 U142 ( .B1(n1050), .B2(n1052), .A(n964), .ZN(n966) );
  INV_X1 U143 ( .A(n966), .ZN(n965) );
  OAI22_X1 U144 ( .A1(A[23]), .A2(n965), .B1(A[23]), .B2(B[28]), .ZN(n967) );
  OAI22_X1 U145 ( .A1(n941), .A2(n967), .B1(n967), .B2(n966), .ZN(n974) );
  OAI221_X1 U146 ( .B1(B[25]), .B2(n968), .C1(A[27]), .C2(B[25]), .A(n974), 
        .ZN(n970) );
  OAI21_X1 U147 ( .B1(A[24]), .B2(A[27]), .A(n940), .ZN(n969) );
  NAND2_X1 U148 ( .A1(A[25]), .A2(B[27]), .ZN(n1020) );
  NAND2_X1 U149 ( .A1(A[26]), .A2(B[26]), .ZN(n1017) );
  AND2_X1 U150 ( .A1(n1020), .A2(n1017), .ZN(n976) );
  NAND3_X1 U151 ( .A1(n970), .A2(n969), .A3(n976), .ZN(n1024) );
  XOR2_X1 U152 ( .A(n1024), .B(n940), .Z(n972) );
  XOR2_X1 U153 ( .A(n941), .B(n1024), .Z(n971) );
  OAI22_X1 U154 ( .A1(n1077), .A2(n972), .B1(A[28]), .B2(n971), .ZN(SUM[28])
         );
  INV_X1 U155 ( .A(n974), .ZN(n1007) );
  OAI21_X1 U156 ( .B1(n1007), .B2(n941), .A(n1076), .ZN(n973) );
  OAI21_X1 U157 ( .B1(B[23]), .B2(n974), .A(n973), .ZN(n1022) );
  INV_X1 U158 ( .A(n975), .ZN(n1016) );
  INV_X1 U159 ( .A(n1015), .ZN(n1021) );
  NAND2_X1 U160 ( .A1(n1016), .A2(n1021), .ZN(n977) );
  OAI21_X1 U161 ( .B1(n1022), .B2(n977), .A(n976), .ZN(n1002) );
  XOR2_X1 U162 ( .A(A[27]), .B(n940), .Z(n978) );
  XOR2_X1 U163 ( .A(n1002), .B(n978), .Z(SUM[27]) );
  XOR2_X1 U164 ( .A(A[24]), .B(n941), .Z(n1008) );
  XOR2_X1 U165 ( .A(n1008), .B(n1007), .Z(SUM[24]) );
  NAND2_X1 U166 ( .A1(n1040), .A2(n1009), .ZN(n1010) );
  XOR2_X1 U167 ( .A(n1010), .B(n940), .Z(n1012) );
  XOR2_X1 U168 ( .A(n941), .B(n1010), .Z(n1011) );
  OAI22_X1 U169 ( .A1(n947), .A2(n1012), .B1(A[19]), .B2(n1011), .ZN(SUM[19])
         );
  OAI21_X1 U170 ( .B1(n1015), .B2(n1022), .A(n1020), .ZN(n1019) );
  AND2_X1 U171 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U172 ( .A(n1019), .B(n1018), .Z(SUM[26]) );
  NAND2_X1 U173 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XOR2_X1 U174 ( .A(n1023), .B(n1022), .Z(SUM[25]) );
  INV_X1 U175 ( .A(A[29]), .ZN(n1026) );
  OAI222_X1 U176 ( .A1(A[28]), .A2(n1024), .B1(A[28]), .B2(B[24]), .C1(B[24]), 
        .C2(n1024), .ZN(n1045) );
  AND2_X1 U177 ( .A1(n1026), .A2(n1045), .ZN(n1025) );
  OAI22_X1 U178 ( .A1(n1026), .A2(n1045), .B1(n1025), .B2(n1041), .ZN(n1032)
         );
  INV_X1 U185 ( .A(n1032), .ZN(n1028) );
  OAI22_X1 U186 ( .A1(A[30]), .A2(B[21]), .B1(n940), .B2(n1032), .ZN(n1027) );
  OAI22_X1 U187 ( .A1(n1028), .A2(n1027), .B1(n1117), .B2(n1027), .ZN(n1030)
         );
  XOR2_X1 U188 ( .A(A[31]), .B(n940), .Z(n1029) );
  XOR2_X1 U189 ( .A(n1030), .B(n1029), .Z(SUM[31]) );
  XOR2_X1 U190 ( .A(A[30]), .B(n940), .Z(n1031) );
  XOR2_X1 U191 ( .A(n1032), .B(n1031), .Z(SUM[30]) );
  NOR2_X1 U192 ( .A1(n1034), .A2(n1033), .ZN(n1037) );
  XOR2_X1 U193 ( .A(n1035), .B(n941), .Z(n1036) );
  XOR2_X1 U194 ( .A(n1037), .B(n1036), .Z(SUM[21]) );
  INV_X1 U195 ( .A(n1038), .ZN(n1039) );
  NAND2_X1 U196 ( .A1(n1040), .A2(n1039), .ZN(n1069) );
  XOR2_X1 U197 ( .A(A[17]), .B(n1041), .Z(n1043) );
  XNOR2_X1 U198 ( .A(n1043), .B(n1042), .ZN(SUM[17]) );
  XOR2_X1 U199 ( .A(B[17]), .B(A[29]), .Z(n1044) );
  XNOR2_X1 U200 ( .A(n1045), .B(n1044), .ZN(SUM[29]) );
  INV_X1 U201 ( .A(n1046), .ZN(n1047) );
  NOR2_X1 U202 ( .A1(n1048), .A2(n1047), .ZN(n1075) );
  NOR2_X1 U203 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XOR2_X1 U204 ( .A(n1052), .B(n1051), .Z(SUM[22]) );
endmodule


module BRANCHDECISIONUNIT ( OPCODE, JOFFSET_IN, BOFFSET_IN, NPC_IN, REG1_IN, 
        REG2_IN, NPC_OUT );
  input [5:0] OPCODE;
  input [25:0] JOFFSET_IN;
  input [15:0] BOFFSET_IN;
  input [31:0] NPC_IN;
  input [31:0] REG1_IN;
  input [31:0] REG2_IN;
  output [31:0] NPC_OUT;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N429, N428, N425, N424, N412, N411, N410, N409, N408,
         N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397,
         N395, N388, N380, N379, N378, N377, N376, N375, N374, N373, N372,
         N371, N370, N369, N368, N367, N366, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443;
  wire   [31:0] boffsetadjusted;
  wire   [31:0] joffsetadjusted;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10;

  NAND3_X1 U178 ( .A1(OPCODE[2]), .A2(n98), .A3(n99), .ZN(n95) );
  NAND3_X1 U179 ( .A1(n98), .A2(n442), .A3(OPCODE[1]), .ZN(n96) );
  BOFFSET BOFF ( .BOFFSET_IN(BOFFSET_IN), .BOFFSET_OUT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, boffsetadjusted[27], 
        SYNOPSYS_UNCONNECTED__4, boffsetadjusted[25:24], 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, boffsetadjusted[20], SYNOPSYS_UNCONNECTED__8, 
        boffsetadjusted[18:17], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, boffsetadjusted[14:0]}) );
  JOFFSET JOFF ( .JOFFSET_IN(JOFFSET_IN), .JOFFSET_OUT(joffsetadjusted) );
  BRANCHDECISIONUNIT_DW01_add_5 r62 ( .A(NPC_IN), .B(joffsetadjusted), .CI(
        1'b0), .SUM({N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, N15, N14, N13, N12}) );
  BRANCHDECISIONUNIT_DW01_add_7 add_59_aco ( .A(NPC_IN), .B({N429, N428, N428, 
        N428, N425, N424, N428, N424, N428, N424, N424, N429, N428, N425, N429, 
        N429, N429, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, 
        N402, N401, N400, N399, N398}), .CI(1'b0), .SUM({N114, N113, N112, 
        N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, 
        N85, N84, N83}) );
  BRANCHDECISIONUNIT_DW01_add_6 add_53_aco ( .A(NPC_IN), .B({n423, n423, N395, 
        n423, n423, n423, n423, n423, n423, N388, n423, N388, n423, n423, N395, 
        N388, N395, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, 
        N370, N369, N368, N367, N366}), .CI(1'b0), .SUM({N78, N77, N76, N75, 
        N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47})
         );
  NAND2_X1 U1 ( .A1(n101), .A2(n102), .ZN(n100) );
  NOR2_X1 U2 ( .A1(n443), .A2(n424), .ZN(N429) );
  AND2_X1 U3 ( .A1(boffsetadjusted[17]), .A2(n443), .ZN(N395) );
  AND2_X1 U7 ( .A1(boffsetadjusted[18]), .A2(n443), .ZN(N388) );
  BUF_X1 U8 ( .A(n30), .Z(n417) );
  BUF_X1 U9 ( .A(n30), .Z(n418) );
  BUF_X1 U10 ( .A(n29), .Z(n420) );
  BUF_X1 U11 ( .A(n29), .Z(n421) );
  BUF_X1 U12 ( .A(n441), .Z(n411) );
  BUF_X1 U13 ( .A(n441), .Z(n412) );
  BUF_X1 U14 ( .A(n440), .Z(n408) );
  BUF_X1 U15 ( .A(n440), .Z(n409) );
  BUF_X1 U16 ( .A(n30), .Z(n419) );
  BUF_X1 U17 ( .A(n29), .Z(n422) );
  BUF_X1 U18 ( .A(n441), .Z(n413) );
  BUF_X1 U19 ( .A(n440), .Z(n410) );
  INV_X1 U20 ( .A(n100), .ZN(n443) );
  NOR2_X1 U21 ( .A1(n443), .A2(n426), .ZN(N399) );
  NOR2_X1 U22 ( .A1(n443), .A2(n428), .ZN(N401) );
  NOR2_X1 U23 ( .A1(n443), .A2(n427), .ZN(N400) );
  NOR2_X1 U24 ( .A1(n443), .A2(n425), .ZN(N398) );
  NOR2_X1 U25 ( .A1(n443), .A2(n436), .ZN(N409) );
  NOR2_X1 U26 ( .A1(n443), .A2(n438), .ZN(N411) );
  NOR2_X1 U27 ( .A1(n443), .A2(n430), .ZN(N403) );
  NOR2_X1 U28 ( .A1(n443), .A2(n434), .ZN(N407) );
  NOR2_X1 U29 ( .A1(n443), .A2(n435), .ZN(N408) );
  NOR2_X1 U30 ( .A1(n443), .A2(n439), .ZN(N412) );
  NOR2_X1 U31 ( .A1(n443), .A2(n437), .ZN(N410) );
  NOR2_X1 U32 ( .A1(n443), .A2(n431), .ZN(N404) );
  NOR2_X1 U33 ( .A1(n443), .A2(n429), .ZN(N402) );
  NOR2_X1 U34 ( .A1(n443), .A2(n432), .ZN(N405) );
  NOR2_X1 U35 ( .A1(n443), .A2(n433), .ZN(N406) );
  NOR2_X1 U36 ( .A1(n427), .A2(n100), .ZN(N368) );
  AND2_X1 U37 ( .A1(boffsetadjusted[25]), .A2(n100), .ZN(N428) );
  NOR2_X1 U38 ( .A1(n430), .A2(n100), .ZN(N371) );
  NOR2_X1 U39 ( .A1(n435), .A2(n100), .ZN(N376) );
  NOR2_X1 U40 ( .A1(n434), .A2(n100), .ZN(N375) );
  NOR2_X1 U41 ( .A1(n433), .A2(n100), .ZN(N374) );
  NOR2_X1 U42 ( .A1(n432), .A2(n100), .ZN(N373) );
  AND2_X1 U43 ( .A1(boffsetadjusted[24]), .A2(n100), .ZN(N424) );
  NOR2_X1 U44 ( .A1(n428), .A2(n100), .ZN(N369) );
  NOR2_X1 U45 ( .A1(n429), .A2(n100), .ZN(N370) );
  NOR2_X1 U46 ( .A1(n431), .A2(n100), .ZN(N372) );
  NOR2_X1 U47 ( .A1(n439), .A2(n100), .ZN(N380) );
  NOR2_X1 U48 ( .A1(n438), .A2(n100), .ZN(N379) );
  NOR2_X1 U49 ( .A1(n425), .A2(n100), .ZN(N366) );
  NOR2_X1 U50 ( .A1(n426), .A2(n100), .ZN(N367) );
  NOR2_X1 U51 ( .A1(n437), .A2(n100), .ZN(N378) );
  AND2_X1 U52 ( .A1(boffsetadjusted[27]), .A2(n100), .ZN(N425) );
  NOR2_X1 U53 ( .A1(n436), .A2(n100), .ZN(N377) );
  BUF_X1 U54 ( .A(N397), .Z(n423) );
  NOR2_X1 U55 ( .A1(n424), .A2(n100), .ZN(N397) );
  NOR2_X1 U56 ( .A1(n96), .A2(n416), .ZN(n30) );
  BUF_X1 U57 ( .A(n31), .Z(n416) );
  BUF_X1 U58 ( .A(n31), .Z(n415) );
  BUF_X1 U59 ( .A(n31), .Z(n414) );
  AND3_X1 U60 ( .A1(n95), .A2(n96), .A3(n94), .ZN(n29) );
  INV_X1 U61 ( .A(n95), .ZN(n440) );
  INV_X1 U62 ( .A(n94), .ZN(n441) );
  NAND2_X1 U63 ( .A1(n54), .A2(n55), .ZN(NPC_OUT[27]) );
  AOI22_X1 U64 ( .A1(REG1_IN[27]), .A2(n418), .B1(N39), .B2(n415), .ZN(n54) );
  AOI222_X1 U65 ( .A1(N74), .A2(n409), .B1(NPC_IN[27]), .B2(n421), .C1(N110), 
        .C2(n412), .ZN(n55) );
  NAND2_X1 U66 ( .A1(n52), .A2(n53), .ZN(NPC_OUT[28]) );
  AOI22_X1 U67 ( .A1(REG1_IN[28]), .A2(n418), .B1(N40), .B2(n414), .ZN(n52) );
  AOI222_X1 U68 ( .A1(N75), .A2(n409), .B1(NPC_IN[28]), .B2(n421), .C1(N111), 
        .C2(n412), .ZN(n53) );
  NAND2_X1 U69 ( .A1(n50), .A2(n51), .ZN(NPC_OUT[29]) );
  AOI22_X1 U70 ( .A1(REG1_IN[29]), .A2(n418), .B1(N41), .B2(n414), .ZN(n50) );
  AOI222_X1 U71 ( .A1(N76), .A2(n409), .B1(NPC_IN[29]), .B2(n421), .C1(N112), 
        .C2(n412), .ZN(n51) );
  NAND2_X1 U72 ( .A1(n46), .A2(n47), .ZN(NPC_OUT[30]) );
  AOI22_X1 U73 ( .A1(REG1_IN[30]), .A2(n418), .B1(N42), .B2(n414), .ZN(n46) );
  AOI222_X1 U74 ( .A1(N77), .A2(n409), .B1(NPC_IN[30]), .B2(n421), .C1(N113), 
        .C2(n412), .ZN(n47) );
  NOR4_X1 U75 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(n102) );
  NOR4_X1 U76 ( .A1(n107), .A2(n108), .A3(n109), .A4(n110), .ZN(n101) );
  OR4_X1 U77 ( .A1(REG1_IN[6]), .A2(REG1_IN[7]), .A3(REG1_IN[8]), .A4(
        REG1_IN[9]), .ZN(n103) );
  NAND2_X1 U78 ( .A1(n44), .A2(n45), .ZN(NPC_OUT[31]) );
  AOI22_X1 U79 ( .A1(REG1_IN[31]), .A2(n419), .B1(N43), .B2(n414), .ZN(n44) );
  AOI222_X1 U80 ( .A1(N78), .A2(n410), .B1(NPC_IN[31]), .B2(n422), .C1(N114), 
        .C2(n413), .ZN(n45) );
  OR4_X1 U81 ( .A1(REG1_IN[0]), .A2(REG1_IN[10]), .A3(REG1_IN[11]), .A4(
        REG1_IN[12]), .ZN(n110) );
  OR4_X1 U82 ( .A1(REG1_IN[24]), .A2(REG1_IN[25]), .A3(REG1_IN[26]), .A4(
        REG1_IN[27]), .ZN(n106) );
  OR4_X1 U83 ( .A1(REG1_IN[13]), .A2(REG1_IN[14]), .A3(REG1_IN[15]), .A4(
        REG1_IN[16]), .ZN(n109) );
  OR4_X1 U84 ( .A1(REG1_IN[28]), .A2(REG1_IN[29]), .A3(REG1_IN[2]), .A4(
        REG1_IN[30]), .ZN(n105) );
  OR4_X1 U85 ( .A1(REG1_IN[17]), .A2(REG1_IN[18]), .A3(REG1_IN[19]), .A4(
        REG1_IN[1]), .ZN(n108) );
  OR4_X1 U86 ( .A1(REG1_IN[31]), .A2(REG1_IN[3]), .A3(REG1_IN[4]), .A4(
        REG1_IN[5]), .ZN(n104) );
  OR4_X1 U87 ( .A1(REG1_IN[20]), .A2(REG1_IN[21]), .A3(REG1_IN[22]), .A4(
        REG1_IN[23]), .ZN(n107) );
  NAND2_X1 U88 ( .A1(n68), .A2(n69), .ZN(NPC_OUT[20]) );
  AOI22_X1 U89 ( .A1(REG1_IN[20]), .A2(n418), .B1(N32), .B2(n415), .ZN(n68) );
  AOI222_X1 U90 ( .A1(N67), .A2(n409), .B1(NPC_IN[20]), .B2(n421), .C1(N103), 
        .C2(n412), .ZN(n69) );
  NAND2_X1 U91 ( .A1(n66), .A2(n67), .ZN(NPC_OUT[21]) );
  AOI22_X1 U92 ( .A1(REG1_IN[21]), .A2(n418), .B1(N33), .B2(n415), .ZN(n66) );
  AOI222_X1 U93 ( .A1(N68), .A2(n409), .B1(NPC_IN[21]), .B2(n421), .C1(N104), 
        .C2(n412), .ZN(n67) );
  NAND2_X1 U94 ( .A1(n64), .A2(n65), .ZN(NPC_OUT[22]) );
  AOI22_X1 U95 ( .A1(REG1_IN[22]), .A2(n418), .B1(N34), .B2(n415), .ZN(n64) );
  AOI222_X1 U96 ( .A1(N69), .A2(n409), .B1(NPC_IN[22]), .B2(n421), .C1(N105), 
        .C2(n412), .ZN(n65) );
  NAND2_X1 U97 ( .A1(n60), .A2(n61), .ZN(NPC_OUT[24]) );
  AOI22_X1 U98 ( .A1(REG1_IN[24]), .A2(n418), .B1(N36), .B2(n415), .ZN(n60) );
  AOI222_X1 U99 ( .A1(N71), .A2(n409), .B1(NPC_IN[24]), .B2(n421), .C1(N107), 
        .C2(n412), .ZN(n61) );
  NAND2_X1 U100 ( .A1(n58), .A2(n59), .ZN(NPC_OUT[25]) );
  AOI22_X1 U101 ( .A1(REG1_IN[25]), .A2(n418), .B1(N37), .B2(n415), .ZN(n58)
         );
  AOI222_X1 U102 ( .A1(N72), .A2(n409), .B1(NPC_IN[25]), .B2(n421), .C1(N108), 
        .C2(n412), .ZN(n59) );
  NAND2_X1 U103 ( .A1(n56), .A2(n57), .ZN(NPC_OUT[26]) );
  AOI22_X1 U104 ( .A1(REG1_IN[26]), .A2(n418), .B1(N38), .B2(n415), .ZN(n56)
         );
  AOI222_X1 U105 ( .A1(N73), .A2(n409), .B1(NPC_IN[26]), .B2(n421), .C1(N109), 
        .C2(n412), .ZN(n57) );
  NAND2_X1 U106 ( .A1(n62), .A2(n63), .ZN(NPC_OUT[23]) );
  AOI22_X1 U107 ( .A1(REG1_IN[23]), .A2(n418), .B1(N35), .B2(n415), .ZN(n62)
         );
  AOI222_X1 U108 ( .A1(N70), .A2(n409), .B1(NPC_IN[23]), .B2(n421), .C1(N106), 
        .C2(n412), .ZN(n63) );
  NAND2_X1 U109 ( .A1(n90), .A2(n91), .ZN(NPC_OUT[10]) );
  AOI22_X1 U110 ( .A1(REG1_IN[10]), .A2(n417), .B1(N22), .B2(n416), .ZN(n90)
         );
  AOI222_X1 U111 ( .A1(N57), .A2(n408), .B1(NPC_IN[10]), .B2(n420), .C1(N93), 
        .C2(n411), .ZN(n91) );
  NAND2_X1 U112 ( .A1(n84), .A2(n85), .ZN(NPC_OUT[13]) );
  AOI22_X1 U113 ( .A1(REG1_IN[13]), .A2(n417), .B1(N25), .B2(n416), .ZN(n84)
         );
  AOI222_X1 U114 ( .A1(N60), .A2(n408), .B1(NPC_IN[13]), .B2(n420), .C1(N96), 
        .C2(n411), .ZN(n85) );
  NAND2_X1 U115 ( .A1(n82), .A2(n83), .ZN(NPC_OUT[14]) );
  AOI22_X1 U116 ( .A1(REG1_IN[14]), .A2(n417), .B1(N26), .B2(n416), .ZN(n82)
         );
  AOI222_X1 U117 ( .A1(N61), .A2(n408), .B1(NPC_IN[14]), .B2(n420), .C1(N97), 
        .C2(n411), .ZN(n83) );
  NAND2_X1 U118 ( .A1(n80), .A2(n81), .ZN(NPC_OUT[15]) );
  AOI22_X1 U119 ( .A1(REG1_IN[15]), .A2(n417), .B1(N27), .B2(n416), .ZN(n80)
         );
  AOI222_X1 U120 ( .A1(N62), .A2(n408), .B1(NPC_IN[15]), .B2(n420), .C1(N98), 
        .C2(n411), .ZN(n81) );
  NAND2_X1 U121 ( .A1(n78), .A2(n79), .ZN(NPC_OUT[16]) );
  AOI22_X1 U122 ( .A1(REG1_IN[16]), .A2(n417), .B1(N28), .B2(n416), .ZN(n78)
         );
  AOI222_X1 U123 ( .A1(N63), .A2(n408), .B1(NPC_IN[16]), .B2(n420), .C1(N99), 
        .C2(n411), .ZN(n79) );
  NAND2_X1 U124 ( .A1(n74), .A2(n75), .ZN(NPC_OUT[18]) );
  AOI22_X1 U125 ( .A1(REG1_IN[18]), .A2(n417), .B1(N30), .B2(n415), .ZN(n74)
         );
  AOI222_X1 U126 ( .A1(N65), .A2(n408), .B1(NPC_IN[18]), .B2(n420), .C1(N101), 
        .C2(n411), .ZN(n75) );
  NAND2_X1 U127 ( .A1(n72), .A2(n73), .ZN(NPC_OUT[19]) );
  AOI22_X1 U128 ( .A1(REG1_IN[19]), .A2(n417), .B1(N31), .B2(n415), .ZN(n72)
         );
  AOI222_X1 U129 ( .A1(N66), .A2(n408), .B1(NPC_IN[19]), .B2(n420), .C1(N102), 
        .C2(n411), .ZN(n73) );
  NAND2_X1 U130 ( .A1(n27), .A2(n28), .ZN(NPC_OUT[9]) );
  AOI22_X1 U131 ( .A1(REG1_IN[9]), .A2(n419), .B1(N21), .B2(n414), .ZN(n27) );
  AOI222_X1 U132 ( .A1(N56), .A2(n410), .B1(NPC_IN[9]), .B2(n422), .C1(N92), 
        .C2(n413), .ZN(n28) );
  NAND2_X1 U133 ( .A1(n76), .A2(n77), .ZN(NPC_OUT[17]) );
  AOI22_X1 U134 ( .A1(REG1_IN[17]), .A2(n417), .B1(N29), .B2(n415), .ZN(n76)
         );
  AOI222_X1 U135 ( .A1(N64), .A2(n408), .B1(NPC_IN[17]), .B2(n420), .C1(N100), 
        .C2(n411), .ZN(n77) );
  NAND2_X1 U136 ( .A1(n32), .A2(n33), .ZN(NPC_OUT[8]) );
  AOI22_X1 U137 ( .A1(REG1_IN[8]), .A2(n419), .B1(N20), .B2(n414), .ZN(n32) );
  AOI222_X1 U138 ( .A1(N55), .A2(n410), .B1(NPC_IN[8]), .B2(n422), .C1(N91), 
        .C2(n413), .ZN(n33) );
  NAND2_X1 U139 ( .A1(n34), .A2(n35), .ZN(NPC_OUT[7]) );
  AOI22_X1 U140 ( .A1(REG1_IN[7]), .A2(n419), .B1(N19), .B2(n414), .ZN(n34) );
  AOI222_X1 U141 ( .A1(N54), .A2(n410), .B1(NPC_IN[7]), .B2(n422), .C1(N90), 
        .C2(n413), .ZN(n35) );
  NAND2_X1 U142 ( .A1(n88), .A2(n89), .ZN(NPC_OUT[11]) );
  AOI22_X1 U143 ( .A1(REG1_IN[11]), .A2(n417), .B1(N23), .B2(n416), .ZN(n88)
         );
  AOI222_X1 U144 ( .A1(N58), .A2(n408), .B1(NPC_IN[11]), .B2(n420), .C1(N94), 
        .C2(n411), .ZN(n89) );
  NAND2_X1 U145 ( .A1(n86), .A2(n87), .ZN(NPC_OUT[12]) );
  AOI22_X1 U146 ( .A1(REG1_IN[12]), .A2(n417), .B1(N24), .B2(n416), .ZN(n86)
         );
  AOI222_X1 U147 ( .A1(N59), .A2(n408), .B1(NPC_IN[12]), .B2(n420), .C1(N95), 
        .C2(n411), .ZN(n87) );
  INV_X1 U148 ( .A(boffsetadjusted[4]), .ZN(n429) );
  INV_X1 U149 ( .A(boffsetadjusted[5]), .ZN(n430) );
  INV_X1 U150 ( .A(boffsetadjusted[6]), .ZN(n431) );
  INV_X1 U151 ( .A(boffsetadjusted[9]), .ZN(n434) );
  INV_X1 U152 ( .A(boffsetadjusted[10]), .ZN(n435) );
  INV_X1 U153 ( .A(boffsetadjusted[8]), .ZN(n433) );
  INV_X1 U154 ( .A(boffsetadjusted[3]), .ZN(n428) );
  INV_X1 U155 ( .A(boffsetadjusted[0]), .ZN(n425) );
  INV_X1 U156 ( .A(boffsetadjusted[1]), .ZN(n426) );
  INV_X1 U157 ( .A(boffsetadjusted[2]), .ZN(n427) );
  NAND2_X1 U158 ( .A1(n38), .A2(n39), .ZN(NPC_OUT[5]) );
  AOI22_X1 U159 ( .A1(REG1_IN[5]), .A2(n419), .B1(N17), .B2(n414), .ZN(n38) );
  AOI222_X1 U160 ( .A1(N52), .A2(n410), .B1(NPC_IN[5]), .B2(n422), .C1(N88), 
        .C2(n413), .ZN(n39) );
  NAND2_X1 U161 ( .A1(n36), .A2(n37), .ZN(NPC_OUT[6]) );
  AOI22_X1 U162 ( .A1(REG1_IN[6]), .A2(n419), .B1(N18), .B2(n414), .ZN(n36) );
  AOI222_X1 U163 ( .A1(N53), .A2(n410), .B1(NPC_IN[6]), .B2(n422), .C1(N89), 
        .C2(n413), .ZN(n37) );
  NAND2_X1 U164 ( .A1(n40), .A2(n41), .ZN(NPC_OUT[4]) );
  AOI22_X1 U165 ( .A1(REG1_IN[4]), .A2(n419), .B1(N16), .B2(n414), .ZN(n40) );
  AOI222_X1 U166 ( .A1(N51), .A2(n410), .B1(NPC_IN[4]), .B2(n422), .C1(N87), 
        .C2(n413), .ZN(n41) );
  NAND2_X1 U167 ( .A1(n48), .A2(n49), .ZN(NPC_OUT[2]) );
  AOI22_X1 U168 ( .A1(REG1_IN[2]), .A2(n418), .B1(N14), .B2(n414), .ZN(n48) );
  AOI222_X1 U169 ( .A1(N49), .A2(n409), .B1(NPC_IN[2]), .B2(n421), .C1(N85), 
        .C2(n412), .ZN(n49) );
  NAND2_X1 U170 ( .A1(n42), .A2(n43), .ZN(NPC_OUT[3]) );
  AOI22_X1 U171 ( .A1(REG1_IN[3]), .A2(n419), .B1(N15), .B2(n414), .ZN(n42) );
  AOI222_X1 U172 ( .A1(N50), .A2(n410), .B1(NPC_IN[3]), .B2(n422), .C1(N86), 
        .C2(n413), .ZN(n43) );
  INV_X1 U173 ( .A(boffsetadjusted[11]), .ZN(n436) );
  INV_X1 U174 ( .A(boffsetadjusted[12]), .ZN(n437) );
  INV_X1 U175 ( .A(boffsetadjusted[13]), .ZN(n438) );
  INV_X1 U176 ( .A(boffsetadjusted[14]), .ZN(n439) );
  INV_X1 U177 ( .A(boffsetadjusted[7]), .ZN(n432) );
  NAND2_X1 U180 ( .A1(n92), .A2(n93), .ZN(NPC_OUT[0]) );
  AOI22_X1 U181 ( .A1(REG1_IN[0]), .A2(n417), .B1(N12), .B2(n416), .ZN(n92) );
  AOI222_X1 U182 ( .A1(N47), .A2(n408), .B1(NPC_IN[0]), .B2(n420), .C1(N83), 
        .C2(n411), .ZN(n93) );
  NAND2_X1 U183 ( .A1(n70), .A2(n71), .ZN(NPC_OUT[1]) );
  AOI22_X1 U184 ( .A1(REG1_IN[1]), .A2(n417), .B1(N13), .B2(n415), .ZN(n70) );
  AOI222_X1 U185 ( .A1(N48), .A2(n408), .B1(NPC_IN[1]), .B2(n420), .C1(N84), 
        .C2(n411), .ZN(n71) );
  INV_X1 U186 ( .A(OPCODE[2]), .ZN(n442) );
  NOR2_X1 U187 ( .A1(n96), .A2(OPCODE[4]), .ZN(n31) );
  NOR2_X1 U188 ( .A1(OPCODE[5]), .A2(OPCODE[3]), .ZN(n98) );
  NOR3_X1 U189 ( .A1(OPCODE[0]), .A2(OPCODE[4]), .A3(OPCODE[1]), .ZN(n99) );
  NAND4_X1 U190 ( .A1(OPCODE[0]), .A2(OPCODE[2]), .A3(n97), .A4(n98), .ZN(n94)
         );
  NOR2_X1 U191 ( .A1(OPCODE[4]), .A2(OPCODE[1]), .ZN(n97) );
  INV_X1 U192 ( .A(boffsetadjusted[20]), .ZN(n424) );
endmodule


module DECODE_STAGE_numbit32 ( IR_IN, WB_STAGE_IN, NPC_IN, RD_IN, CLK, RESET, 
        WRITE_ENABLE, INSTRUCTION_FETCHED, NPC_OUT_BPU, RD_OUT, NPC_OUT, 
        A_REG_OUT, B_REG_OUT, IMM_REG_OUT, alu_forwarding_one, 
        mem_forwarding_one, alu_forwarding_two, mem_forwarding_two );
  input [31:0] IR_IN;
  input [31:0] WB_STAGE_IN;
  input [31:0] NPC_IN;
  input [4:0] RD_IN;
  input [31:0] INSTRUCTION_FETCHED;
  output [31:0] NPC_OUT_BPU;
  output [4:0] RD_OUT;
  output [31:0] NPC_OUT;
  output [31:0] A_REG_OUT;
  output [31:0] B_REG_OUT;
  output [31:0] IMM_REG_OUT;
  input CLK, RESET, WRITE_ENABLE;
  output alu_forwarding_one, mem_forwarding_one, alu_forwarding_two,
         mem_forwarding_two;
  wire   n76, n77;
  wire   [31:0] sign_extention_signal;
  wire   [31:0] RF_ONE_OUT;
  wire   [31:0] RF_TWO_OUT;
  wire   [4:0] rdmux_out;

  SIGN_EXTENTION SIGN_REG ( .D({n76, IR_IN[14:0]}), .Q(sign_extention_signal)
         );
  REGISTER_FILE_numBit_data32_numBit_address5_numBit_registers32 RF ( .CK(CLK), 
        .Reset(n77), .Write_enable(WRITE_ENABLE), .Write_address(RD_IN), 
        .Read_one_address(IR_IN[25:21]), .Read_two_address(IR_IN[20:16]), 
        .Data_in(WB_STAGE_IN), .Data_one_out(RF_ONE_OUT), .Data_two_out(
        RF_TWO_OUT) );
  REGISTER_GENERIC_NBIT32_7 REGONE ( .D(RF_ONE_OUT), .CK(CLK), .RESET(n77), 
        .Q(A_REG_OUT) );
  REGISTER_GENERIC_NBIT32_6 REGTWO ( .D(RF_TWO_OUT), .CK(CLK), .RESET(n77), 
        .Q(B_REG_OUT) );
  REGISTER_GENERIC_NBIT32_5 IMMREG ( .D(sign_extention_signal), .CK(CLK), 
        .RESET(n77), .Q(IMM_REG_OUT) );
  REGISTER_GENERIC_NBIT32_4 NPC_REG ( .D(NPC_IN), .CK(CLK), .RESET(n77), .Q(
        NPC_OUT) );
  RDMUX RDMUX_MUX ( .rtype_in({n76, IR_IN[14:11]}), .itype_in(IR_IN[20:16]), 
        .opcode_in(IR_IN[31:26]), .rd_out(rdmux_out) );
  REGISTER_GENERIC_NBIT5_0 RD_OUT_REG ( .D(rdmux_out), .CK(CLK), .RESET(n77), 
        .Q(RD_OUT) );
  HAZARD_DETECTION HAZARD ( .clk(CLK), .reset(n77), .OPCODE(
        INSTRUCTION_FETCHED[31:26]), .RD_REG_IN_ITYPE(
        INSTRUCTION_FETCHED[20:16]), .RD_REG_IN_RTYPE(
        INSTRUCTION_FETCHED[15:11]), .RS1_REG_IN(INSTRUCTION_FETCHED[25:21]), 
        .RS2_REG_IN(INSTRUCTION_FETCHED[20:16]), .alu_forwarding_one(
        alu_forwarding_one), .mem_forwarding_one(mem_forwarding_one), 
        .alu_forwarding_two(alu_forwarding_two), .mem_forwarding_two(
        mem_forwarding_two) );
  BRANCHDECISIONUNIT BRANCHUNIT ( .OPCODE(IR_IN[31:26]), .JOFFSET_IN({
        IR_IN[25:16], n76, IR_IN[14:0]}), .BOFFSET_IN({n76, IR_IN[14:0]}), 
        .NPC_IN(NPC_IN), .REG1_IN(RF_ONE_OUT), .REG2_IN(RF_TWO_OUT), .NPC_OUT(
        NPC_OUT_BPU) );
  BUF_X1 U1 ( .A(RESET), .Z(n77) );
  BUF_X1 U2 ( .A(IR_IN[15]), .Z(n76) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;

  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_0 UIV_0 ( .A(SEL), .Y(SEL_INV[0]) );
  ND2_0 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_686 UND2_0 ( .A(B[0]), .B(SEL), .Y(NAND_TWO_OUT[0]) );
  ND2_685 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_228 UIV_1 ( .A(SEL), .Y(SEL_INV[1]) );
  ND2_684 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_683 UND2_1 ( .A(B[1]), .B(SEL), .Y(NAND_TWO_OUT[1]) );
  ND2_682 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_227 UIV_2 ( .A(SEL), .Y(SEL_INV[2]) );
  ND2_681 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_680 UND2_2 ( .A(B[2]), .B(SEL), .Y(NAND_TWO_OUT[2]) );
  ND2_679 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_226 UIV_3 ( .A(SEL), .Y(SEL_INV[3]) );
  ND2_678 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_677 UND2_3 ( .A(B[3]), .B(SEL), .Y(NAND_TWO_OUT[3]) );
  ND2_676 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_225 UIV_4 ( .A(SEL), .Y(SEL_INV[4]) );
  ND2_675 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_674 UND2_4 ( .A(B[4]), .B(SEL), .Y(NAND_TWO_OUT[4]) );
  ND2_673 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_224 UIV_5 ( .A(SEL), .Y(SEL_INV[5]) );
  ND2_672 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_671 UND2_5 ( .A(B[5]), .B(SEL), .Y(NAND_TWO_OUT[5]) );
  ND2_670 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_223 UIV_6 ( .A(SEL), .Y(SEL_INV[6]) );
  ND2_669 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_668 UND2_6 ( .A(B[6]), .B(SEL), .Y(NAND_TWO_OUT[6]) );
  ND2_667 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_222 UIV_7 ( .A(SEL), .Y(SEL_INV[7]) );
  ND2_666 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_665 UND2_7 ( .A(B[7]), .B(SEL), .Y(NAND_TWO_OUT[7]) );
  ND2_664 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_221 UIV_8 ( .A(SEL), .Y(SEL_INV[8]) );
  ND2_663 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_662 UND2_8 ( .A(B[8]), .B(SEL), .Y(NAND_TWO_OUT[8]) );
  ND2_661 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_220 UIV_9 ( .A(SEL), .Y(SEL_INV[9]) );
  ND2_660 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_659 UND2_9 ( .A(B[9]), .B(SEL), .Y(NAND_TWO_OUT[9]) );
  ND2_658 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_219 UIV_10 ( .A(SEL), .Y(SEL_INV[10]) );
  ND2_657 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_656 UND2_10 ( .A(B[10]), .B(SEL), .Y(NAND_TWO_OUT[10]) );
  ND2_655 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_218 UIV_11 ( .A(SEL), .Y(SEL_INV[11]) );
  ND2_654 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_653 UND2_11 ( .A(B[11]), .B(SEL), .Y(NAND_TWO_OUT[11]) );
  ND2_652 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_217 UIV_12 ( .A(SEL), .Y(SEL_INV[12]) );
  ND2_651 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_650 UND2_12 ( .A(B[12]), .B(SEL), .Y(NAND_TWO_OUT[12]) );
  ND2_649 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_216 UIV_13 ( .A(SEL), .Y(SEL_INV[13]) );
  ND2_648 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_647 UND2_13 ( .A(B[13]), .B(SEL), .Y(NAND_TWO_OUT[13]) );
  ND2_646 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_215 UIV_14 ( .A(SEL), .Y(SEL_INV[14]) );
  ND2_645 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_644 UND2_14 ( .A(B[14]), .B(SEL), .Y(NAND_TWO_OUT[14]) );
  ND2_643 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_214 UIV_15 ( .A(SEL), .Y(SEL_INV[15]) );
  ND2_642 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_641 UND2_15 ( .A(B[15]), .B(SEL), .Y(NAND_TWO_OUT[15]) );
  ND2_640 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_213 UIV_16 ( .A(SEL), .Y(SEL_INV[16]) );
  ND2_639 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_638 UND2_16 ( .A(B[16]), .B(SEL), .Y(NAND_TWO_OUT[16]) );
  ND2_637 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_212 UIV_17 ( .A(SEL), .Y(SEL_INV[17]) );
  ND2_636 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_635 UND2_17 ( .A(B[17]), .B(SEL), .Y(NAND_TWO_OUT[17]) );
  ND2_634 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_211 UIV_18 ( .A(SEL), .Y(SEL_INV[18]) );
  ND2_633 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_632 UND2_18 ( .A(B[18]), .B(SEL), .Y(NAND_TWO_OUT[18]) );
  ND2_631 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_210 UIV_19 ( .A(SEL), .Y(SEL_INV[19]) );
  ND2_630 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_629 UND2_19 ( .A(B[19]), .B(SEL), .Y(NAND_TWO_OUT[19]) );
  ND2_628 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_209 UIV_20 ( .A(SEL), .Y(SEL_INV[20]) );
  ND2_627 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_626 UND2_20 ( .A(B[20]), .B(SEL), .Y(NAND_TWO_OUT[20]) );
  ND2_625 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_208 UIV_21 ( .A(SEL), .Y(SEL_INV[21]) );
  ND2_624 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_623 UND2_21 ( .A(B[21]), .B(SEL), .Y(NAND_TWO_OUT[21]) );
  ND2_622 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_207 UIV_22 ( .A(SEL), .Y(SEL_INV[22]) );
  ND2_621 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_620 UND2_22 ( .A(B[22]), .B(SEL), .Y(NAND_TWO_OUT[22]) );
  ND2_619 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_206 UIV_23 ( .A(SEL), .Y(SEL_INV[23]) );
  ND2_618 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_617 UND2_23 ( .A(B[23]), .B(SEL), .Y(NAND_TWO_OUT[23]) );
  ND2_616 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_205 UIV_24 ( .A(SEL), .Y(SEL_INV[24]) );
  ND2_615 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_614 UND2_24 ( .A(B[24]), .B(SEL), .Y(NAND_TWO_OUT[24]) );
  ND2_613 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_204 UIV_25 ( .A(SEL), .Y(SEL_INV[25]) );
  ND2_612 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_611 UND2_25 ( .A(B[25]), .B(SEL), .Y(NAND_TWO_OUT[25]) );
  ND2_610 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_203 UIV_26 ( .A(SEL), .Y(SEL_INV[26]) );
  ND2_609 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_608 UND2_26 ( .A(B[26]), .B(SEL), .Y(NAND_TWO_OUT[26]) );
  ND2_607 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_202 UIV_27 ( .A(SEL), .Y(SEL_INV[27]) );
  ND2_606 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_605 UND2_27 ( .A(B[27]), .B(SEL), .Y(NAND_TWO_OUT[27]) );
  ND2_604 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_201 UIV_28 ( .A(SEL), .Y(SEL_INV[28]) );
  ND2_603 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_602 UND2_28 ( .A(B[28]), .B(SEL), .Y(NAND_TWO_OUT[28]) );
  ND2_601 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_200 UIV_29 ( .A(SEL), .Y(SEL_INV[29]) );
  ND2_600 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_599 UND2_29 ( .A(B[29]), .B(SEL), .Y(NAND_TWO_OUT[29]) );
  ND2_598 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_199 UIV_30 ( .A(SEL), .Y(SEL_INV[30]) );
  ND2_597 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_596 UND2_30 ( .A(B[30]), .B(SEL), .Y(NAND_TWO_OUT[30]) );
  ND2_595 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_198 UIV_31 ( .A(SEL), .Y(SEL_INV[31]) );
  ND2_594 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_593 UND2_31 ( .A(B[31]), .B(SEL), .Y(NAND_TWO_OUT[31]) );
  ND2_592 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n43, n44, n45, n46, n47, n48, n49;
  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_197 UIV_0 ( .A(n47), .Y(SEL_INV[0]) );
  ND2_591 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_590 UND2_0 ( .A(B[0]), .B(n45), .Y(NAND_TWO_OUT[0]) );
  ND2_589 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_196 UIV_1 ( .A(n47), .Y(SEL_INV[1]) );
  ND2_588 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_587 UND2_1 ( .A(B[1]), .B(n45), .Y(NAND_TWO_OUT[1]) );
  ND2_586 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_195 UIV_2 ( .A(n47), .Y(SEL_INV[2]) );
  ND2_585 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_584 UND2_2 ( .A(B[2]), .B(n45), .Y(NAND_TWO_OUT[2]) );
  ND2_583 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_194 UIV_3 ( .A(n47), .Y(SEL_INV[3]) );
  ND2_582 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_581 UND2_3 ( .A(B[3]), .B(n45), .Y(NAND_TWO_OUT[3]) );
  ND2_580 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_193 UIV_4 ( .A(n47), .Y(SEL_INV[4]) );
  ND2_579 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_578 UND2_4 ( .A(B[4]), .B(n45), .Y(NAND_TWO_OUT[4]) );
  ND2_577 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_192 UIV_5 ( .A(n47), .Y(SEL_INV[5]) );
  ND2_576 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_575 UND2_5 ( .A(B[5]), .B(n45), .Y(NAND_TWO_OUT[5]) );
  ND2_574 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_191 UIV_6 ( .A(n48), .Y(SEL_INV[6]) );
  ND2_573 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_572 UND2_6 ( .A(B[6]), .B(n45), .Y(NAND_TWO_OUT[6]) );
  ND2_571 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_190 UIV_7 ( .A(n48), .Y(SEL_INV[7]) );
  ND2_570 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_569 UND2_7 ( .A(B[7]), .B(n45), .Y(NAND_TWO_OUT[7]) );
  ND2_568 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_189 UIV_8 ( .A(n48), .Y(SEL_INV[8]) );
  ND2_567 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_566 UND2_8 ( .A(B[8]), .B(n45), .Y(NAND_TWO_OUT[8]) );
  ND2_565 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_188 UIV_9 ( .A(n48), .Y(SEL_INV[9]) );
  ND2_564 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_563 UND2_9 ( .A(B[9]), .B(n45), .Y(NAND_TWO_OUT[9]) );
  ND2_562 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_187 UIV_10 ( .A(n48), .Y(SEL_INV[10]) );
  ND2_561 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_560 UND2_10 ( .A(B[10]), .B(n45), .Y(NAND_TWO_OUT[10]) );
  ND2_559 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_186 UIV_11 ( .A(n48), .Y(SEL_INV[11]) );
  ND2_558 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_557 UND2_11 ( .A(B[11]), .B(n45), .Y(NAND_TWO_OUT[11]) );
  ND2_556 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_185 UIV_12 ( .A(n48), .Y(SEL_INV[12]) );
  ND2_555 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_554 UND2_12 ( .A(B[12]), .B(n46), .Y(NAND_TWO_OUT[12]) );
  ND2_553 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_184 UIV_13 ( .A(n48), .Y(SEL_INV[13]) );
  ND2_552 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_551 UND2_13 ( .A(B[13]), .B(n46), .Y(NAND_TWO_OUT[13]) );
  ND2_550 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_183 UIV_14 ( .A(n48), .Y(SEL_INV[14]) );
  ND2_549 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_548 UND2_14 ( .A(B[14]), .B(n46), .Y(NAND_TWO_OUT[14]) );
  ND2_547 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_182 UIV_15 ( .A(n48), .Y(SEL_INV[15]) );
  ND2_546 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_545 UND2_15 ( .A(B[15]), .B(n46), .Y(NAND_TWO_OUT[15]) );
  ND2_544 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_181 UIV_16 ( .A(n48), .Y(SEL_INV[16]) );
  ND2_543 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_542 UND2_16 ( .A(B[16]), .B(n46), .Y(NAND_TWO_OUT[16]) );
  ND2_541 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_180 UIV_17 ( .A(n48), .Y(SEL_INV[17]) );
  ND2_540 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_539 UND2_17 ( .A(B[17]), .B(n46), .Y(NAND_TWO_OUT[17]) );
  ND2_538 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_179 UIV_18 ( .A(n48), .Y(SEL_INV[18]) );
  ND2_537 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_536 UND2_18 ( .A(B[18]), .B(n46), .Y(NAND_TWO_OUT[18]) );
  ND2_535 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_178 UIV_19 ( .A(n48), .Y(SEL_INV[19]) );
  ND2_534 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_533 UND2_19 ( .A(B[19]), .B(n46), .Y(NAND_TWO_OUT[19]) );
  ND2_532 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_177 UIV_20 ( .A(n48), .Y(SEL_INV[20]) );
  ND2_531 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_530 UND2_20 ( .A(B[20]), .B(n46), .Y(NAND_TWO_OUT[20]) );
  ND2_529 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_176 UIV_21 ( .A(n48), .Y(SEL_INV[21]) );
  ND2_528 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_527 UND2_21 ( .A(B[21]), .B(n46), .Y(NAND_TWO_OUT[21]) );
  ND2_526 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_175 UIV_22 ( .A(n48), .Y(SEL_INV[22]) );
  ND2_525 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_524 UND2_22 ( .A(B[22]), .B(n46), .Y(NAND_TWO_OUT[22]) );
  ND2_523 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_174 UIV_23 ( .A(n49), .Y(SEL_INV[23]) );
  ND2_522 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_521 UND2_23 ( .A(B[23]), .B(n46), .Y(NAND_TWO_OUT[23]) );
  ND2_520 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_173 UIV_24 ( .A(n49), .Y(SEL_INV[24]) );
  ND2_519 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_518 UND2_24 ( .A(B[24]), .B(n47), .Y(NAND_TWO_OUT[24]) );
  ND2_517 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_172 UIV_25 ( .A(n49), .Y(SEL_INV[25]) );
  ND2_516 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_515 UND2_25 ( .A(B[25]), .B(n47), .Y(NAND_TWO_OUT[25]) );
  ND2_514 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_171 UIV_26 ( .A(n49), .Y(SEL_INV[26]) );
  ND2_513 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_512 UND2_26 ( .A(B[26]), .B(n47), .Y(NAND_TWO_OUT[26]) );
  ND2_511 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_170 UIV_27 ( .A(n49), .Y(SEL_INV[27]) );
  ND2_510 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_509 UND2_27 ( .A(B[27]), .B(n47), .Y(NAND_TWO_OUT[27]) );
  ND2_508 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_169 UIV_28 ( .A(n49), .Y(SEL_INV[28]) );
  ND2_507 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_506 UND2_28 ( .A(B[28]), .B(n47), .Y(NAND_TWO_OUT[28]) );
  ND2_505 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_168 UIV_29 ( .A(n49), .Y(SEL_INV[29]) );
  ND2_504 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_503 UND2_29 ( .A(B[29]), .B(n47), .Y(NAND_TWO_OUT[29]) );
  ND2_502 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_167 UIV_30 ( .A(n49), .Y(SEL_INV[30]) );
  ND2_501 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_500 UND2_30 ( .A(B[30]), .B(n47), .Y(NAND_TWO_OUT[30]) );
  ND2_499 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_166 UIV_31 ( .A(n49), .Y(SEL_INV[31]) );
  ND2_498 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_497 UND2_31 ( .A(B[31]), .B(n47), .Y(NAND_TWO_OUT[31]) );
  ND2_496 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n43), .Z(n45) );
  BUF_X1 U2 ( .A(n43), .Z(n46) );
  BUF_X1 U3 ( .A(n43), .Z(n47) );
  BUF_X1 U4 ( .A(n44), .Z(n48) );
  BUF_X1 U5 ( .A(n44), .Z(n49) );
  BUF_X1 U6 ( .A(SEL), .Z(n43) );
  BUF_X1 U7 ( .A(SEL), .Z(n44) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n43, n44, n45, n46, n47, n48, n49;
  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_165 UIV_0 ( .A(n47), .Y(SEL_INV[0]) );
  ND2_495 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_494 UND2_0 ( .A(B[0]), .B(n45), .Y(NAND_TWO_OUT[0]) );
  ND2_493 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_164 UIV_1 ( .A(n47), .Y(SEL_INV[1]) );
  ND2_492 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_491 UND2_1 ( .A(B[1]), .B(n45), .Y(NAND_TWO_OUT[1]) );
  ND2_490 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_163 UIV_2 ( .A(n47), .Y(SEL_INV[2]) );
  ND2_489 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_488 UND2_2 ( .A(B[2]), .B(n45), .Y(NAND_TWO_OUT[2]) );
  ND2_487 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_162 UIV_3 ( .A(n47), .Y(SEL_INV[3]) );
  ND2_486 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_485 UND2_3 ( .A(B[3]), .B(n45), .Y(NAND_TWO_OUT[3]) );
  ND2_484 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_161 UIV_4 ( .A(n47), .Y(SEL_INV[4]) );
  ND2_483 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_482 UND2_4 ( .A(B[4]), .B(n45), .Y(NAND_TWO_OUT[4]) );
  ND2_481 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_160 UIV_5 ( .A(n47), .Y(SEL_INV[5]) );
  ND2_480 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_479 UND2_5 ( .A(B[5]), .B(n45), .Y(NAND_TWO_OUT[5]) );
  ND2_478 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_159 UIV_6 ( .A(n48), .Y(SEL_INV[6]) );
  ND2_477 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_476 UND2_6 ( .A(B[6]), .B(n45), .Y(NAND_TWO_OUT[6]) );
  ND2_475 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_158 UIV_7 ( .A(n48), .Y(SEL_INV[7]) );
  ND2_474 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_473 UND2_7 ( .A(B[7]), .B(n45), .Y(NAND_TWO_OUT[7]) );
  ND2_472 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_157 UIV_8 ( .A(n48), .Y(SEL_INV[8]) );
  ND2_471 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_470 UND2_8 ( .A(B[8]), .B(n45), .Y(NAND_TWO_OUT[8]) );
  ND2_469 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_156 UIV_9 ( .A(n48), .Y(SEL_INV[9]) );
  ND2_468 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_467 UND2_9 ( .A(B[9]), .B(n45), .Y(NAND_TWO_OUT[9]) );
  ND2_466 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_155 UIV_10 ( .A(n48), .Y(SEL_INV[10]) );
  ND2_465 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_464 UND2_10 ( .A(B[10]), .B(n45), .Y(NAND_TWO_OUT[10]) );
  ND2_463 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_154 UIV_11 ( .A(n48), .Y(SEL_INV[11]) );
  ND2_462 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_461 UND2_11 ( .A(B[11]), .B(n45), .Y(NAND_TWO_OUT[11]) );
  ND2_460 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_153 UIV_12 ( .A(n48), .Y(SEL_INV[12]) );
  ND2_459 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_458 UND2_12 ( .A(B[12]), .B(n46), .Y(NAND_TWO_OUT[12]) );
  ND2_457 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_152 UIV_13 ( .A(n48), .Y(SEL_INV[13]) );
  ND2_456 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_455 UND2_13 ( .A(B[13]), .B(n46), .Y(NAND_TWO_OUT[13]) );
  ND2_454 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_151 UIV_14 ( .A(n48), .Y(SEL_INV[14]) );
  ND2_453 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_452 UND2_14 ( .A(B[14]), .B(n46), .Y(NAND_TWO_OUT[14]) );
  ND2_451 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_150 UIV_15 ( .A(n48), .Y(SEL_INV[15]) );
  ND2_450 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_449 UND2_15 ( .A(B[15]), .B(n46), .Y(NAND_TWO_OUT[15]) );
  ND2_448 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_149 UIV_16 ( .A(n48), .Y(SEL_INV[16]) );
  ND2_447 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_446 UND2_16 ( .A(B[16]), .B(n46), .Y(NAND_TWO_OUT[16]) );
  ND2_445 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_148 UIV_17 ( .A(n48), .Y(SEL_INV[17]) );
  ND2_444 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_443 UND2_17 ( .A(B[17]), .B(n46), .Y(NAND_TWO_OUT[17]) );
  ND2_442 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_147 UIV_18 ( .A(n48), .Y(SEL_INV[18]) );
  ND2_441 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_440 UND2_18 ( .A(B[18]), .B(n46), .Y(NAND_TWO_OUT[18]) );
  ND2_439 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_146 UIV_19 ( .A(n48), .Y(SEL_INV[19]) );
  ND2_438 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_437 UND2_19 ( .A(B[19]), .B(n46), .Y(NAND_TWO_OUT[19]) );
  ND2_436 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_145 UIV_20 ( .A(n48), .Y(SEL_INV[20]) );
  ND2_435 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_434 UND2_20 ( .A(B[20]), .B(n46), .Y(NAND_TWO_OUT[20]) );
  ND2_433 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_144 UIV_21 ( .A(n48), .Y(SEL_INV[21]) );
  ND2_432 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_431 UND2_21 ( .A(B[21]), .B(n46), .Y(NAND_TWO_OUT[21]) );
  ND2_430 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_143 UIV_22 ( .A(n48), .Y(SEL_INV[22]) );
  ND2_429 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_428 UND2_22 ( .A(B[22]), .B(n46), .Y(NAND_TWO_OUT[22]) );
  ND2_427 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_142 UIV_23 ( .A(n49), .Y(SEL_INV[23]) );
  ND2_426 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_425 UND2_23 ( .A(B[23]), .B(n46), .Y(NAND_TWO_OUT[23]) );
  ND2_424 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_141 UIV_24 ( .A(n49), .Y(SEL_INV[24]) );
  ND2_423 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_422 UND2_24 ( .A(B[24]), .B(n47), .Y(NAND_TWO_OUT[24]) );
  ND2_421 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_140 UIV_25 ( .A(n49), .Y(SEL_INV[25]) );
  ND2_420 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_419 UND2_25 ( .A(B[25]), .B(n47), .Y(NAND_TWO_OUT[25]) );
  ND2_418 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_139 UIV_26 ( .A(n49), .Y(SEL_INV[26]) );
  ND2_417 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_416 UND2_26 ( .A(B[26]), .B(n47), .Y(NAND_TWO_OUT[26]) );
  ND2_415 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_138 UIV_27 ( .A(n49), .Y(SEL_INV[27]) );
  ND2_414 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_413 UND2_27 ( .A(B[27]), .B(n47), .Y(NAND_TWO_OUT[27]) );
  ND2_412 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_137 UIV_28 ( .A(n49), .Y(SEL_INV[28]) );
  ND2_411 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_410 UND2_28 ( .A(B[28]), .B(n47), .Y(NAND_TWO_OUT[28]) );
  ND2_409 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_136 UIV_29 ( .A(n49), .Y(SEL_INV[29]) );
  ND2_408 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_407 UND2_29 ( .A(B[29]), .B(n47), .Y(NAND_TWO_OUT[29]) );
  ND2_406 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_135 UIV_30 ( .A(n49), .Y(SEL_INV[30]) );
  ND2_405 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_404 UND2_30 ( .A(B[30]), .B(n47), .Y(NAND_TWO_OUT[30]) );
  ND2_403 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_134 UIV_31 ( .A(n49), .Y(SEL_INV[31]) );
  ND2_402 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_401 UND2_31 ( .A(B[31]), .B(n47), .Y(NAND_TWO_OUT[31]) );
  ND2_400 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n43), .Z(n45) );
  BUF_X1 U2 ( .A(n43), .Z(n46) );
  BUF_X1 U3 ( .A(n43), .Z(n47) );
  BUF_X1 U4 ( .A(n44), .Z(n48) );
  BUF_X1 U5 ( .A(n44), .Z(n49) );
  BUF_X1 U6 ( .A(SEL), .Z(n43) );
  BUF_X1 U7 ( .A(SEL), .Z(n44) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;

  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_133 UIV_0 ( .A(SEL), .Y(SEL_INV[0]) );
  ND2_399 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_398 UND2_0 ( .A(B[0]), .B(SEL), .Y(NAND_TWO_OUT[0]) );
  ND2_397 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_132 UIV_1 ( .A(SEL), .Y(SEL_INV[1]) );
  ND2_396 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_395 UND2_1 ( .A(B[1]), .B(SEL), .Y(NAND_TWO_OUT[1]) );
  ND2_394 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_131 UIV_2 ( .A(SEL), .Y(SEL_INV[2]) );
  ND2_393 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_392 UND2_2 ( .A(B[2]), .B(SEL), .Y(NAND_TWO_OUT[2]) );
  ND2_391 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_130 UIV_3 ( .A(SEL), .Y(SEL_INV[3]) );
  ND2_390 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_389 UND2_3 ( .A(B[3]), .B(SEL), .Y(NAND_TWO_OUT[3]) );
  ND2_388 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_129 UIV_4 ( .A(SEL), .Y(SEL_INV[4]) );
  ND2_387 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_386 UND2_4 ( .A(B[4]), .B(SEL), .Y(NAND_TWO_OUT[4]) );
  ND2_385 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_128 UIV_5 ( .A(SEL), .Y(SEL_INV[5]) );
  ND2_384 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_383 UND2_5 ( .A(B[5]), .B(SEL), .Y(NAND_TWO_OUT[5]) );
  ND2_382 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_127 UIV_6 ( .A(SEL), .Y(SEL_INV[6]) );
  ND2_381 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_380 UND2_6 ( .A(B[6]), .B(SEL), .Y(NAND_TWO_OUT[6]) );
  ND2_379 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_126 UIV_7 ( .A(SEL), .Y(SEL_INV[7]) );
  ND2_378 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_377 UND2_7 ( .A(B[7]), .B(SEL), .Y(NAND_TWO_OUT[7]) );
  ND2_376 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_125 UIV_8 ( .A(SEL), .Y(SEL_INV[8]) );
  ND2_375 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_374 UND2_8 ( .A(B[8]), .B(SEL), .Y(NAND_TWO_OUT[8]) );
  ND2_373 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_124 UIV_9 ( .A(SEL), .Y(SEL_INV[9]) );
  ND2_372 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_371 UND2_9 ( .A(B[9]), .B(SEL), .Y(NAND_TWO_OUT[9]) );
  ND2_370 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_123 UIV_10 ( .A(SEL), .Y(SEL_INV[10]) );
  ND2_369 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_368 UND2_10 ( .A(B[10]), .B(SEL), .Y(NAND_TWO_OUT[10]) );
  ND2_367 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_122 UIV_11 ( .A(SEL), .Y(SEL_INV[11]) );
  ND2_366 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_365 UND2_11 ( .A(B[11]), .B(SEL), .Y(NAND_TWO_OUT[11]) );
  ND2_364 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_121 UIV_12 ( .A(SEL), .Y(SEL_INV[12]) );
  ND2_363 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_362 UND2_12 ( .A(B[12]), .B(SEL), .Y(NAND_TWO_OUT[12]) );
  ND2_361 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_120 UIV_13 ( .A(SEL), .Y(SEL_INV[13]) );
  ND2_360 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_359 UND2_13 ( .A(B[13]), .B(SEL), .Y(NAND_TWO_OUT[13]) );
  ND2_358 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_119 UIV_14 ( .A(SEL), .Y(SEL_INV[14]) );
  ND2_357 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_356 UND2_14 ( .A(B[14]), .B(SEL), .Y(NAND_TWO_OUT[14]) );
  ND2_355 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_118 UIV_15 ( .A(SEL), .Y(SEL_INV[15]) );
  ND2_354 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_353 UND2_15 ( .A(B[15]), .B(SEL), .Y(NAND_TWO_OUT[15]) );
  ND2_352 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_117 UIV_16 ( .A(SEL), .Y(SEL_INV[16]) );
  ND2_351 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_350 UND2_16 ( .A(B[16]), .B(SEL), .Y(NAND_TWO_OUT[16]) );
  ND2_349 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_116 UIV_17 ( .A(SEL), .Y(SEL_INV[17]) );
  ND2_348 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_347 UND2_17 ( .A(B[17]), .B(SEL), .Y(NAND_TWO_OUT[17]) );
  ND2_346 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_115 UIV_18 ( .A(SEL), .Y(SEL_INV[18]) );
  ND2_345 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_344 UND2_18 ( .A(B[18]), .B(SEL), .Y(NAND_TWO_OUT[18]) );
  ND2_343 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_114 UIV_19 ( .A(SEL), .Y(SEL_INV[19]) );
  ND2_342 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_341 UND2_19 ( .A(B[19]), .B(SEL), .Y(NAND_TWO_OUT[19]) );
  ND2_340 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_113 UIV_20 ( .A(SEL), .Y(SEL_INV[20]) );
  ND2_339 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_338 UND2_20 ( .A(B[20]), .B(SEL), .Y(NAND_TWO_OUT[20]) );
  ND2_337 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_112 UIV_21 ( .A(SEL), .Y(SEL_INV[21]) );
  ND2_336 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_335 UND2_21 ( .A(B[21]), .B(SEL), .Y(NAND_TWO_OUT[21]) );
  ND2_334 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_111 UIV_22 ( .A(SEL), .Y(SEL_INV[22]) );
  ND2_333 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_332 UND2_22 ( .A(B[22]), .B(SEL), .Y(NAND_TWO_OUT[22]) );
  ND2_331 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_110 UIV_23 ( .A(SEL), .Y(SEL_INV[23]) );
  ND2_330 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_329 UND2_23 ( .A(B[23]), .B(SEL), .Y(NAND_TWO_OUT[23]) );
  ND2_328 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_109 UIV_24 ( .A(SEL), .Y(SEL_INV[24]) );
  ND2_327 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_326 UND2_24 ( .A(B[24]), .B(SEL), .Y(NAND_TWO_OUT[24]) );
  ND2_325 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_108 UIV_25 ( .A(SEL), .Y(SEL_INV[25]) );
  ND2_324 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_323 UND2_25 ( .A(B[25]), .B(SEL), .Y(NAND_TWO_OUT[25]) );
  ND2_322 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_107 UIV_26 ( .A(SEL), .Y(SEL_INV[26]) );
  ND2_321 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_320 UND2_26 ( .A(B[26]), .B(SEL), .Y(NAND_TWO_OUT[26]) );
  ND2_319 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_106 UIV_27 ( .A(SEL), .Y(SEL_INV[27]) );
  ND2_318 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_317 UND2_27 ( .A(B[27]), .B(SEL), .Y(NAND_TWO_OUT[27]) );
  ND2_316 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_105 UIV_28 ( .A(SEL), .Y(SEL_INV[28]) );
  ND2_315 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_314 UND2_28 ( .A(B[28]), .B(SEL), .Y(NAND_TWO_OUT[28]) );
  ND2_313 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_104 UIV_29 ( .A(SEL), .Y(SEL_INV[29]) );
  ND2_312 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_311 UND2_29 ( .A(B[29]), .B(SEL), .Y(NAND_TWO_OUT[29]) );
  ND2_310 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_103 UIV_30 ( .A(SEL), .Y(SEL_INV[30]) );
  ND2_309 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_308 UND2_30 ( .A(B[30]), .B(SEL), .Y(NAND_TWO_OUT[30]) );
  ND2_307 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_102 UIV_31 ( .A(SEL), .Y(SEL_INV[31]) );
  ND2_306 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_305 UND2_31 ( .A(B[31]), .B(SEL), .Y(NAND_TWO_OUT[31]) );
  ND2_304 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n43, n44, n45, n46, n47, n48, n49;
  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_101 UIV_0 ( .A(n47), .Y(SEL_INV[0]) );
  ND2_303 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_302 UND2_0 ( .A(B[0]), .B(n45), .Y(NAND_TWO_OUT[0]) );
  ND2_301 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_100 UIV_1 ( .A(n47), .Y(SEL_INV[1]) );
  ND2_300 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_299 UND2_1 ( .A(B[1]), .B(n45), .Y(NAND_TWO_OUT[1]) );
  ND2_298 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_99 UIV_2 ( .A(n47), .Y(SEL_INV[2]) );
  ND2_297 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_296 UND2_2 ( .A(B[2]), .B(n45), .Y(NAND_TWO_OUT[2]) );
  ND2_295 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_98 UIV_3 ( .A(n47), .Y(SEL_INV[3]) );
  ND2_294 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_293 UND2_3 ( .A(B[3]), .B(n45), .Y(NAND_TWO_OUT[3]) );
  ND2_292 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_97 UIV_4 ( .A(n47), .Y(SEL_INV[4]) );
  ND2_291 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_290 UND2_4 ( .A(B[4]), .B(n45), .Y(NAND_TWO_OUT[4]) );
  ND2_289 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_96 UIV_5 ( .A(n47), .Y(SEL_INV[5]) );
  ND2_288 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_287 UND2_5 ( .A(B[5]), .B(n45), .Y(NAND_TWO_OUT[5]) );
  ND2_286 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_95 UIV_6 ( .A(n48), .Y(SEL_INV[6]) );
  ND2_285 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_284 UND2_6 ( .A(B[6]), .B(n45), .Y(NAND_TWO_OUT[6]) );
  ND2_283 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_94 UIV_7 ( .A(n48), .Y(SEL_INV[7]) );
  ND2_282 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_281 UND2_7 ( .A(B[7]), .B(n45), .Y(NAND_TWO_OUT[7]) );
  ND2_280 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_93 UIV_8 ( .A(n48), .Y(SEL_INV[8]) );
  ND2_279 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_278 UND2_8 ( .A(B[8]), .B(n45), .Y(NAND_TWO_OUT[8]) );
  ND2_277 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_92 UIV_9 ( .A(n48), .Y(SEL_INV[9]) );
  ND2_276 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_275 UND2_9 ( .A(B[9]), .B(n45), .Y(NAND_TWO_OUT[9]) );
  ND2_274 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_91 UIV_10 ( .A(n48), .Y(SEL_INV[10]) );
  ND2_273 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_272 UND2_10 ( .A(B[10]), .B(n45), .Y(NAND_TWO_OUT[10]) );
  ND2_271 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_90 UIV_11 ( .A(n48), .Y(SEL_INV[11]) );
  ND2_270 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_269 UND2_11 ( .A(B[11]), .B(n45), .Y(NAND_TWO_OUT[11]) );
  ND2_268 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_89 UIV_12 ( .A(n48), .Y(SEL_INV[12]) );
  ND2_267 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_266 UND2_12 ( .A(B[12]), .B(n46), .Y(NAND_TWO_OUT[12]) );
  ND2_265 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_88 UIV_13 ( .A(n48), .Y(SEL_INV[13]) );
  ND2_264 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_263 UND2_13 ( .A(B[13]), .B(n46), .Y(NAND_TWO_OUT[13]) );
  ND2_262 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_87 UIV_14 ( .A(n48), .Y(SEL_INV[14]) );
  ND2_261 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_260 UND2_14 ( .A(B[14]), .B(n46), .Y(NAND_TWO_OUT[14]) );
  ND2_259 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_86 UIV_15 ( .A(n48), .Y(SEL_INV[15]) );
  ND2_258 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_257 UND2_15 ( .A(B[15]), .B(n46), .Y(NAND_TWO_OUT[15]) );
  ND2_256 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_85 UIV_16 ( .A(n48), .Y(SEL_INV[16]) );
  ND2_255 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_254 UND2_16 ( .A(B[16]), .B(n46), .Y(NAND_TWO_OUT[16]) );
  ND2_253 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_84 UIV_17 ( .A(n48), .Y(SEL_INV[17]) );
  ND2_252 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_251 UND2_17 ( .A(B[17]), .B(n46), .Y(NAND_TWO_OUT[17]) );
  ND2_250 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_83 UIV_18 ( .A(n48), .Y(SEL_INV[18]) );
  ND2_249 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_248 UND2_18 ( .A(B[18]), .B(n46), .Y(NAND_TWO_OUT[18]) );
  ND2_247 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_82 UIV_19 ( .A(n48), .Y(SEL_INV[19]) );
  ND2_246 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_245 UND2_19 ( .A(B[19]), .B(n46), .Y(NAND_TWO_OUT[19]) );
  ND2_244 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_81 UIV_20 ( .A(n48), .Y(SEL_INV[20]) );
  ND2_243 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_242 UND2_20 ( .A(B[20]), .B(n46), .Y(NAND_TWO_OUT[20]) );
  ND2_241 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_80 UIV_21 ( .A(n48), .Y(SEL_INV[21]) );
  ND2_240 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_239 UND2_21 ( .A(B[21]), .B(n46), .Y(NAND_TWO_OUT[21]) );
  ND2_238 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_79 UIV_22 ( .A(n48), .Y(SEL_INV[22]) );
  ND2_237 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_236 UND2_22 ( .A(B[22]), .B(n46), .Y(NAND_TWO_OUT[22]) );
  ND2_235 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_78 UIV_23 ( .A(n49), .Y(SEL_INV[23]) );
  ND2_234 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_233 UND2_23 ( .A(B[23]), .B(n46), .Y(NAND_TWO_OUT[23]) );
  ND2_232 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_77 UIV_24 ( .A(n49), .Y(SEL_INV[24]) );
  ND2_231 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_230 UND2_24 ( .A(B[24]), .B(n47), .Y(NAND_TWO_OUT[24]) );
  ND2_229 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_76 UIV_25 ( .A(n49), .Y(SEL_INV[25]) );
  ND2_228 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_227 UND2_25 ( .A(B[25]), .B(n47), .Y(NAND_TWO_OUT[25]) );
  ND2_226 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_75 UIV_26 ( .A(n49), .Y(SEL_INV[26]) );
  ND2_225 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_224 UND2_26 ( .A(B[26]), .B(n47), .Y(NAND_TWO_OUT[26]) );
  ND2_223 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_74 UIV_27 ( .A(n49), .Y(SEL_INV[27]) );
  ND2_222 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_221 UND2_27 ( .A(B[27]), .B(n47), .Y(NAND_TWO_OUT[27]) );
  ND2_220 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_73 UIV_28 ( .A(n49), .Y(SEL_INV[28]) );
  ND2_219 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_218 UND2_28 ( .A(B[28]), .B(n47), .Y(NAND_TWO_OUT[28]) );
  ND2_217 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_72 UIV_29 ( .A(n49), .Y(SEL_INV[29]) );
  ND2_216 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_215 UND2_29 ( .A(B[29]), .B(n47), .Y(NAND_TWO_OUT[29]) );
  ND2_214 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_71 UIV_30 ( .A(n49), .Y(SEL_INV[30]) );
  ND2_213 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_212 UND2_30 ( .A(B[30]), .B(n47), .Y(NAND_TWO_OUT[30]) );
  ND2_211 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_70 UIV_31 ( .A(n49), .Y(SEL_INV[31]) );
  ND2_210 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_209 UND2_31 ( .A(B[31]), .B(n47), .Y(NAND_TWO_OUT[31]) );
  ND2_208 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n43), .Z(n45) );
  BUF_X1 U2 ( .A(n43), .Z(n47) );
  BUF_X1 U3 ( .A(n43), .Z(n46) );
  BUF_X1 U4 ( .A(n44), .Z(n48) );
  BUF_X1 U5 ( .A(n44), .Z(n49) );
  BUF_X1 U6 ( .A(SEL), .Z(n43) );
  BUF_X1 U7 ( .A(SEL), .Z(n44) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n43, n44, n45, n46, n47, n48, n49;
  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_69 UIV_0 ( .A(n47), .Y(SEL_INV[0]) );
  ND2_207 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_206 UND2_0 ( .A(B[0]), .B(n45), .Y(NAND_TWO_OUT[0]) );
  ND2_205 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_68 UIV_1 ( .A(n47), .Y(SEL_INV[1]) );
  ND2_204 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_203 UND2_1 ( .A(B[1]), .B(n45), .Y(NAND_TWO_OUT[1]) );
  ND2_202 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_67 UIV_2 ( .A(n47), .Y(SEL_INV[2]) );
  ND2_201 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_200 UND2_2 ( .A(B[2]), .B(n45), .Y(NAND_TWO_OUT[2]) );
  ND2_199 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_66 UIV_3 ( .A(n47), .Y(SEL_INV[3]) );
  ND2_198 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_197 UND2_3 ( .A(B[3]), .B(n45), .Y(NAND_TWO_OUT[3]) );
  ND2_196 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_65 UIV_4 ( .A(n47), .Y(SEL_INV[4]) );
  ND2_195 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_194 UND2_4 ( .A(B[4]), .B(n45), .Y(NAND_TWO_OUT[4]) );
  ND2_193 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_64 UIV_5 ( .A(n47), .Y(SEL_INV[5]) );
  ND2_192 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_191 UND2_5 ( .A(B[5]), .B(n45), .Y(NAND_TWO_OUT[5]) );
  ND2_190 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_63 UIV_6 ( .A(n48), .Y(SEL_INV[6]) );
  ND2_189 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_188 UND2_6 ( .A(B[6]), .B(n45), .Y(NAND_TWO_OUT[6]) );
  ND2_187 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_62 UIV_7 ( .A(n48), .Y(SEL_INV[7]) );
  ND2_186 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_185 UND2_7 ( .A(B[7]), .B(n45), .Y(NAND_TWO_OUT[7]) );
  ND2_184 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_61 UIV_8 ( .A(n48), .Y(SEL_INV[8]) );
  ND2_183 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_182 UND2_8 ( .A(B[8]), .B(n45), .Y(NAND_TWO_OUT[8]) );
  ND2_181 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_60 UIV_9 ( .A(n48), .Y(SEL_INV[9]) );
  ND2_180 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_179 UND2_9 ( .A(B[9]), .B(n45), .Y(NAND_TWO_OUT[9]) );
  ND2_178 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_59 UIV_10 ( .A(n48), .Y(SEL_INV[10]) );
  ND2_177 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_176 UND2_10 ( .A(B[10]), .B(n45), .Y(NAND_TWO_OUT[10]) );
  ND2_175 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_58 UIV_11 ( .A(n48), .Y(SEL_INV[11]) );
  ND2_174 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_173 UND2_11 ( .A(B[11]), .B(n45), .Y(NAND_TWO_OUT[11]) );
  ND2_172 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_57 UIV_12 ( .A(n48), .Y(SEL_INV[12]) );
  ND2_171 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_170 UND2_12 ( .A(B[12]), .B(n46), .Y(NAND_TWO_OUT[12]) );
  ND2_169 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_56 UIV_13 ( .A(n48), .Y(SEL_INV[13]) );
  ND2_168 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_167 UND2_13 ( .A(B[13]), .B(n46), .Y(NAND_TWO_OUT[13]) );
  ND2_166 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_55 UIV_14 ( .A(n48), .Y(SEL_INV[14]) );
  ND2_165 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_164 UND2_14 ( .A(B[14]), .B(n46), .Y(NAND_TWO_OUT[14]) );
  ND2_163 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_54 UIV_15 ( .A(n48), .Y(SEL_INV[15]) );
  ND2_162 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_161 UND2_15 ( .A(B[15]), .B(n46), .Y(NAND_TWO_OUT[15]) );
  ND2_160 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_53 UIV_16 ( .A(n48), .Y(SEL_INV[16]) );
  ND2_159 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_158 UND2_16 ( .A(B[16]), .B(n46), .Y(NAND_TWO_OUT[16]) );
  ND2_157 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_52 UIV_17 ( .A(n48), .Y(SEL_INV[17]) );
  ND2_156 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_155 UND2_17 ( .A(B[17]), .B(n46), .Y(NAND_TWO_OUT[17]) );
  ND2_154 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_51 UIV_18 ( .A(n48), .Y(SEL_INV[18]) );
  ND2_153 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_152 UND2_18 ( .A(B[18]), .B(n46), .Y(NAND_TWO_OUT[18]) );
  ND2_151 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_50 UIV_19 ( .A(n48), .Y(SEL_INV[19]) );
  ND2_150 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_149 UND2_19 ( .A(B[19]), .B(n46), .Y(NAND_TWO_OUT[19]) );
  ND2_148 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_49 UIV_20 ( .A(n48), .Y(SEL_INV[20]) );
  ND2_147 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_146 UND2_20 ( .A(B[20]), .B(n46), .Y(NAND_TWO_OUT[20]) );
  ND2_145 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_48 UIV_21 ( .A(n48), .Y(SEL_INV[21]) );
  ND2_144 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_143 UND2_21 ( .A(B[21]), .B(n46), .Y(NAND_TWO_OUT[21]) );
  ND2_142 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_47 UIV_22 ( .A(n48), .Y(SEL_INV[22]) );
  ND2_141 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_140 UND2_22 ( .A(B[22]), .B(n46), .Y(NAND_TWO_OUT[22]) );
  ND2_139 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_46 UIV_23 ( .A(n49), .Y(SEL_INV[23]) );
  ND2_138 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_137 UND2_23 ( .A(B[23]), .B(n46), .Y(NAND_TWO_OUT[23]) );
  ND2_136 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_45 UIV_24 ( .A(n49), .Y(SEL_INV[24]) );
  ND2_135 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_134 UND2_24 ( .A(B[24]), .B(n47), .Y(NAND_TWO_OUT[24]) );
  ND2_133 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_44 UIV_25 ( .A(n49), .Y(SEL_INV[25]) );
  ND2_132 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_131 UND2_25 ( .A(B[25]), .B(n47), .Y(NAND_TWO_OUT[25]) );
  ND2_130 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_43 UIV_26 ( .A(n49), .Y(SEL_INV[26]) );
  ND2_129 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_128 UND2_26 ( .A(B[26]), .B(n47), .Y(NAND_TWO_OUT[26]) );
  ND2_127 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_42 UIV_27 ( .A(n49), .Y(SEL_INV[27]) );
  ND2_126 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_125 UND2_27 ( .A(B[27]), .B(n47), .Y(NAND_TWO_OUT[27]) );
  ND2_124 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_41 UIV_28 ( .A(n49), .Y(SEL_INV[28]) );
  ND2_123 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_122 UND2_28 ( .A(B[28]), .B(n47), .Y(NAND_TWO_OUT[28]) );
  ND2_121 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_40 UIV_29 ( .A(n49), .Y(SEL_INV[29]) );
  ND2_120 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_119 UND2_29 ( .A(B[29]), .B(n47), .Y(NAND_TWO_OUT[29]) );
  ND2_118 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_39 UIV_30 ( .A(n49), .Y(SEL_INV[30]) );
  ND2_117 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_116 UND2_30 ( .A(B[30]), .B(n47), .Y(NAND_TWO_OUT[30]) );
  ND2_115 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_38 UIV_31 ( .A(n49), .Y(SEL_INV[31]) );
  ND2_114 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_113 UND2_31 ( .A(B[31]), .B(n47), .Y(NAND_TWO_OUT[31]) );
  ND2_112 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n43), .Z(n45) );
  BUF_X1 U2 ( .A(n43), .Z(n47) );
  BUF_X1 U3 ( .A(n43), .Z(n46) );
  BUF_X1 U4 ( .A(n44), .Z(n48) );
  BUF_X1 U5 ( .A(n44), .Z(n49) );
  BUF_X1 U6 ( .A(SEL), .Z(n43) );
  BUF_X1 U7 ( .A(SEL), .Z(n44) );
endmodule


module ALU_BEHAVIORAL_NBIT32_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226;
  wire   [32:0] carry;

  FA_X1 U2_31 ( .A(A[31]), .B(n226), .CI(carry[31]), .S(DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n225), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n224), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n223), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n222), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n221), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n220), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n219), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n218), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n217), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n216), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n215), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n214), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n213), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n212), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n211), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n210), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n209), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n208), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n207), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n206), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n205), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n204), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n203), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FA_X1 U2_7 ( .A(A[7]), .B(n202), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FA_X1 U2_6 ( .A(A[6]), .B(n201), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FA_X1 U2_5 ( .A(A[5]), .B(n200), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FA_X1 U2_4 ( .A(A[4]), .B(n199), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FA_X1 U2_3 ( .A(A[3]), .B(n198), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FA_X1 U2_2 ( .A(A[2]), .B(n197), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FA_X1 U2_1 ( .A(A[1]), .B(n196), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(DIFF[0]) );
  INV_X1 U2 ( .A(B[1]), .ZN(n196) );
  NAND2_X1 U3 ( .A1(B[0]), .A2(n195), .ZN(carry[1]) );
  INV_X1 U4 ( .A(A[0]), .ZN(n195) );
  INV_X1 U5 ( .A(B[2]), .ZN(n197) );
  INV_X1 U6 ( .A(B[3]), .ZN(n198) );
  INV_X1 U7 ( .A(B[4]), .ZN(n199) );
  INV_X1 U8 ( .A(B[5]), .ZN(n200) );
  INV_X1 U9 ( .A(B[6]), .ZN(n201) );
  INV_X1 U10 ( .A(B[7]), .ZN(n202) );
  INV_X1 U11 ( .A(B[8]), .ZN(n203) );
  INV_X1 U12 ( .A(B[9]), .ZN(n204) );
  INV_X1 U13 ( .A(B[10]), .ZN(n205) );
  INV_X1 U14 ( .A(B[11]), .ZN(n206) );
  INV_X1 U15 ( .A(B[12]), .ZN(n207) );
  INV_X1 U16 ( .A(B[13]), .ZN(n208) );
  INV_X1 U17 ( .A(B[14]), .ZN(n209) );
  INV_X1 U18 ( .A(B[15]), .ZN(n210) );
  INV_X1 U19 ( .A(B[16]), .ZN(n211) );
  INV_X1 U20 ( .A(B[17]), .ZN(n212) );
  INV_X1 U21 ( .A(B[18]), .ZN(n213) );
  INV_X1 U22 ( .A(B[19]), .ZN(n214) );
  INV_X1 U23 ( .A(B[20]), .ZN(n215) );
  INV_X1 U24 ( .A(B[21]), .ZN(n216) );
  INV_X1 U25 ( .A(B[22]), .ZN(n217) );
  INV_X1 U26 ( .A(B[23]), .ZN(n218) );
  INV_X1 U27 ( .A(B[24]), .ZN(n219) );
  INV_X1 U28 ( .A(B[25]), .ZN(n220) );
  INV_X1 U29 ( .A(B[26]), .ZN(n221) );
  INV_X1 U30 ( .A(B[27]), .ZN(n222) );
  INV_X1 U31 ( .A(B[28]), .ZN(n223) );
  INV_X1 U32 ( .A(B[29]), .ZN(n224) );
  INV_X1 U33 ( .A(B[30]), .ZN(n225) );
  INV_X1 U34 ( .A(B[31]), .ZN(n226) );
endmodule


module ALU_BEHAVIORAL_NBIT32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
endmodule


module ALU_BEHAVIORAL_NBIT32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n530, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XOR2_X1 U103 ( .A(A[30]), .B(n591), .Z(n70) );
  NAND3_X1 U172 ( .A1(n197), .A2(n150), .A3(n147), .ZN(n196) );
  NAND3_X1 U176 ( .A1(n536), .A2(n199), .A3(n200), .ZN(n197) );
  INV_X1 U1 ( .A(n130), .ZN(n549) );
  INV_X1 U2 ( .A(n118), .ZN(n557) );
  INV_X1 U3 ( .A(n106), .ZN(n565) );
  INV_X1 U4 ( .A(n94), .ZN(n573) );
  INV_X1 U5 ( .A(n82), .ZN(n581) );
  INV_X1 U6 ( .A(n142), .ZN(n541) );
  NOR2_X1 U7 ( .A1(n193), .A2(n136), .ZN(n135) );
  NOR2_X1 U8 ( .A1(n187), .A2(n124), .ZN(n123) );
  NOR2_X1 U9 ( .A1(n181), .A2(n112), .ZN(n111) );
  NOR2_X1 U10 ( .A1(n175), .A2(n100), .ZN(n99) );
  NOR2_X1 U11 ( .A1(n169), .A2(n88), .ZN(n87) );
  NOR2_X1 U12 ( .A1(n163), .A2(n76), .ZN(n75) );
  OAI211_X1 U13 ( .C1(n161), .C2(n162), .A(n78), .B(n75), .ZN(n160) );
  NAND2_X1 U14 ( .A1(n584), .A2(n164), .ZN(n162) );
  AOI211_X1 U15 ( .C1(n165), .C2(n166), .A(n82), .B(n579), .ZN(n161) );
  INV_X1 U16 ( .A(n79), .ZN(n584) );
  OAI211_X1 U17 ( .C1(n191), .C2(n192), .A(n138), .B(n135), .ZN(n190) );
  NAND2_X1 U18 ( .A1(n544), .A2(n194), .ZN(n192) );
  AOI211_X1 U19 ( .C1(n195), .C2(n196), .A(n142), .B(n539), .ZN(n191) );
  INV_X1 U20 ( .A(n139), .ZN(n544) );
  OAI211_X1 U21 ( .C1(n185), .C2(n186), .A(n126), .B(n123), .ZN(n184) );
  NAND2_X1 U22 ( .A1(n552), .A2(n188), .ZN(n186) );
  AOI211_X1 U23 ( .C1(n189), .C2(n190), .A(n130), .B(n547), .ZN(n185) );
  INV_X1 U24 ( .A(n127), .ZN(n552) );
  OAI211_X1 U25 ( .C1(n179), .C2(n180), .A(n114), .B(n111), .ZN(n178) );
  NAND2_X1 U26 ( .A1(n560), .A2(n182), .ZN(n180) );
  AOI211_X1 U27 ( .C1(n183), .C2(n184), .A(n118), .B(n555), .ZN(n179) );
  INV_X1 U28 ( .A(n115), .ZN(n560) );
  OAI211_X1 U29 ( .C1(n173), .C2(n174), .A(n102), .B(n99), .ZN(n172) );
  NAND2_X1 U30 ( .A1(n568), .A2(n176), .ZN(n174) );
  AOI211_X1 U31 ( .C1(n177), .C2(n178), .A(n106), .B(n563), .ZN(n173) );
  INV_X1 U32 ( .A(n103), .ZN(n568) );
  OAI211_X1 U33 ( .C1(n167), .C2(n168), .A(n90), .B(n87), .ZN(n166) );
  NAND2_X1 U34 ( .A1(n576), .A2(n170), .ZN(n168) );
  AOI211_X1 U35 ( .C1(n171), .C2(n172), .A(n94), .B(n571), .ZN(n167) );
  INV_X1 U36 ( .A(n91), .ZN(n576) );
  AOI21_X1 U37 ( .B1(n143), .B2(n144), .A(n145), .ZN(n140) );
  AOI21_X1 U38 ( .B1(n146), .B2(n147), .A(n148), .ZN(n143) );
  AOI21_X1 U39 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U40 ( .B1(n152), .B2(n153), .A(n534), .ZN(n149) );
  AOI21_X1 U41 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  AOI21_X1 U42 ( .B1(n134), .B2(n135), .A(n136), .ZN(n131) );
  AOI21_X1 U43 ( .B1(n137), .B2(n138), .A(n139), .ZN(n134) );
  AOI21_X1 U44 ( .B1(n140), .B2(n541), .A(n542), .ZN(n137) );
  AOI21_X1 U45 ( .B1(n119), .B2(n120), .A(n121), .ZN(n116) );
  AOI21_X1 U46 ( .B1(n122), .B2(n123), .A(n124), .ZN(n119) );
  AOI21_X1 U47 ( .B1(n125), .B2(n126), .A(n127), .ZN(n122) );
  AOI21_X1 U48 ( .B1(n128), .B2(n549), .A(n550), .ZN(n125) );
  AOI21_X1 U49 ( .B1(n107), .B2(n108), .A(n109), .ZN(n104) );
  AOI21_X1 U50 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  AOI21_X1 U51 ( .B1(n113), .B2(n114), .A(n115), .ZN(n110) );
  AOI21_X1 U52 ( .B1(n116), .B2(n557), .A(n558), .ZN(n113) );
  AOI21_X1 U53 ( .B1(n95), .B2(n96), .A(n97), .ZN(n92) );
  AOI21_X1 U54 ( .B1(n98), .B2(n99), .A(n100), .ZN(n95) );
  AOI21_X1 U55 ( .B1(n101), .B2(n102), .A(n103), .ZN(n98) );
  AOI21_X1 U56 ( .B1(n104), .B2(n565), .A(n566), .ZN(n101) );
  AOI21_X1 U57 ( .B1(n83), .B2(n84), .A(n85), .ZN(n80) );
  AOI21_X1 U58 ( .B1(n86), .B2(n87), .A(n88), .ZN(n83) );
  AOI21_X1 U59 ( .B1(n89), .B2(n90), .A(n91), .ZN(n86) );
  AOI21_X1 U60 ( .B1(n92), .B2(n573), .A(n574), .ZN(n89) );
  AOI21_X1 U61 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI21_X1 U62 ( .B1(n74), .B2(n75), .A(n76), .ZN(n71) );
  AOI21_X1 U63 ( .B1(n77), .B2(n78), .A(n79), .ZN(n74) );
  AOI21_X1 U64 ( .B1(n80), .B2(n581), .A(n582), .ZN(n77) );
  NOR2_X1 U65 ( .A1(n198), .A2(n148), .ZN(n147) );
  NOR2_X1 U66 ( .A1(n198), .A2(n145), .ZN(n195) );
  NOR2_X1 U67 ( .A1(n193), .A2(n133), .ZN(n189) );
  NOR2_X1 U68 ( .A1(n187), .A2(n121), .ZN(n183) );
  NOR2_X1 U69 ( .A1(n181), .A2(n109), .ZN(n177) );
  NOR2_X1 U70 ( .A1(n175), .A2(n97), .ZN(n171) );
  NOR2_X1 U71 ( .A1(n169), .A2(n85), .ZN(n165) );
  NOR2_X1 U72 ( .A1(n163), .A2(n73), .ZN(n159) );
  NAND2_X1 U73 ( .A1(LE), .A2(GE), .ZN(NE) );
  NAND2_X1 U74 ( .A1(n188), .A2(n129), .ZN(n130) );
  NAND2_X1 U75 ( .A1(n182), .A2(n117), .ZN(n118) );
  NAND2_X1 U76 ( .A1(n170), .A2(n93), .ZN(n94) );
  NAND2_X1 U77 ( .A1(n164), .A2(n81), .ZN(n82) );
  NAND2_X1 U78 ( .A1(n176), .A2(n105), .ZN(n106) );
  NAND2_X1 U79 ( .A1(n194), .A2(n141), .ZN(n142) );
  AND2_X1 U80 ( .A1(n199), .A2(n154), .ZN(n153) );
  INV_X1 U81 ( .A(GT), .ZN(LE) );
  INV_X1 U82 ( .A(n132), .ZN(n547) );
  INV_X1 U83 ( .A(n120), .ZN(n555) );
  INV_X1 U84 ( .A(n108), .ZN(n563) );
  INV_X1 U85 ( .A(n96), .ZN(n571) );
  INV_X1 U86 ( .A(n84), .ZN(n579) );
  INV_X1 U87 ( .A(n154), .ZN(n534) );
  INV_X1 U88 ( .A(n144), .ZN(n539) );
  INV_X1 U89 ( .A(n129), .ZN(n550) );
  INV_X1 U90 ( .A(n117), .ZN(n558) );
  INV_X1 U91 ( .A(n93), .ZN(n574) );
  INV_X1 U92 ( .A(n81), .ZN(n582) );
  INV_X1 U93 ( .A(n105), .ZN(n566) );
  INV_X1 U94 ( .A(n141), .ZN(n542) );
  AOI21_X1 U95 ( .B1(n66), .B2(n530), .A(n67), .ZN(GE) );
  INV_X1 U96 ( .A(n68), .ZN(n530) );
  AOI22_X1 U97 ( .A1(B[30]), .A2(n589), .B1(n69), .B2(n70), .ZN(n68) );
  INV_X1 U98 ( .A(A[30]), .ZN(n589) );
  NOR2_X1 U99 ( .A1(n537), .A2(B[3]), .ZN(n151) );
  OAI21_X1 U100 ( .B1(n67), .B2(n157), .A(n66), .ZN(GT) );
  AOI22_X1 U101 ( .A1(A[30]), .A2(n591), .B1(n158), .B2(n70), .ZN(n157) );
  AOI21_X1 U102 ( .B1(n159), .B2(n160), .A(n587), .ZN(n158) );
  INV_X1 U104 ( .A(n72), .ZN(n587) );
  NOR2_X1 U105 ( .A1(n533), .A2(B[0]), .ZN(n201) );
  NOR2_X1 U106 ( .A1(n538), .A2(B[4]), .ZN(n198) );
  NOR2_X1 U107 ( .A1(n592), .A2(A[31]), .ZN(n67) );
  NOR2_X1 U108 ( .A1(n546), .A2(B[8]), .ZN(n193) );
  NOR2_X1 U109 ( .A1(n562), .A2(B[16]), .ZN(n181) );
  NOR2_X1 U110 ( .A1(n578), .A2(B[24]), .ZN(n169) );
  NOR2_X1 U111 ( .A1(n554), .A2(B[12]), .ZN(n187) );
  NOR2_X1 U112 ( .A1(n570), .A2(B[20]), .ZN(n175) );
  NOR2_X1 U113 ( .A1(n586), .A2(B[28]), .ZN(n163) );
  NOR2_X1 U114 ( .A1(n548), .A2(B[9]), .ZN(n133) );
  NOR2_X1 U115 ( .A1(n556), .A2(B[13]), .ZN(n121) );
  NOR2_X1 U116 ( .A1(n564), .A2(B[17]), .ZN(n109) );
  NOR2_X1 U117 ( .A1(n572), .A2(B[21]), .ZN(n97) );
  NOR2_X1 U118 ( .A1(n580), .A2(B[25]), .ZN(n85) );
  AOI22_X1 U119 ( .A1(n155), .A2(n590), .B1(A[1]), .B2(n156), .ZN(n152) );
  OR2_X1 U120 ( .A1(n156), .A2(A[1]), .ZN(n155) );
  NAND2_X1 U121 ( .A1(B[0]), .A2(n533), .ZN(n156) );
  NOR2_X1 U122 ( .A1(n577), .A2(B[23]), .ZN(n91) );
  NOR2_X1 U123 ( .A1(n553), .A2(B[11]), .ZN(n127) );
  NOR2_X1 U124 ( .A1(n585), .A2(B[27]), .ZN(n79) );
  NOR2_X1 U125 ( .A1(n561), .A2(B[15]), .ZN(n115) );
  NOR2_X1 U126 ( .A1(n569), .A2(B[19]), .ZN(n103) );
  NOR2_X1 U127 ( .A1(n540), .A2(B[5]), .ZN(n145) );
  NOR2_X1 U128 ( .A1(n588), .A2(B[29]), .ZN(n73) );
  NOR2_X1 U129 ( .A1(n545), .A2(B[7]), .ZN(n139) );
  NAND2_X1 U130 ( .A1(B[3]), .A2(n537), .ZN(n150) );
  NAND2_X1 U131 ( .A1(A[31]), .A2(n592), .ZN(n66) );
  INV_X1 U132 ( .A(A[3]), .ZN(n537) );
  INV_X1 U133 ( .A(A[11]), .ZN(n553) );
  INV_X1 U134 ( .A(A[27]), .ZN(n585) );
  INV_X1 U135 ( .A(A[9]), .ZN(n548) );
  INV_X1 U136 ( .A(A[13]), .ZN(n556) );
  INV_X1 U137 ( .A(A[17]), .ZN(n564) );
  INV_X1 U138 ( .A(A[21]), .ZN(n572) );
  INV_X1 U139 ( .A(A[23]), .ZN(n577) );
  INV_X1 U140 ( .A(A[25]), .ZN(n580) );
  INV_X1 U141 ( .A(A[15]), .ZN(n561) );
  INV_X1 U142 ( .A(A[19]), .ZN(n569) );
  INV_X1 U143 ( .A(n151), .ZN(n536) );
  OAI211_X1 U144 ( .C1(A[1]), .C2(n201), .A(n532), .B(n153), .ZN(n200) );
  NAND2_X1 U145 ( .A1(B[2]), .A2(n535), .ZN(n154) );
  INV_X1 U146 ( .A(A[5]), .ZN(n540) );
  INV_X1 U147 ( .A(A[7]), .ZN(n545) );
  INV_X1 U148 ( .A(A[26]), .ZN(n583) );
  INV_X1 U149 ( .A(B[1]), .ZN(n590) );
  NAND2_X1 U150 ( .A1(B[23]), .A2(n577), .ZN(n90) );
  NAND2_X1 U151 ( .A1(B[11]), .A2(n553), .ZN(n126) );
  NAND2_X1 U152 ( .A1(B[27]), .A2(n585), .ZN(n78) );
  NAND2_X1 U153 ( .A1(B[15]), .A2(n561), .ZN(n114) );
  NAND2_X1 U154 ( .A1(B[19]), .A2(n569), .ZN(n102) );
  NAND2_X1 U155 ( .A1(B[9]), .A2(n548), .ZN(n132) );
  NAND2_X1 U156 ( .A1(B[13]), .A2(n556), .ZN(n120) );
  NAND2_X1 U157 ( .A1(B[17]), .A2(n564), .ZN(n108) );
  NAND2_X1 U158 ( .A1(B[21]), .A2(n572), .ZN(n96) );
  NAND2_X1 U159 ( .A1(B[25]), .A2(n580), .ZN(n84) );
  INV_X1 U160 ( .A(A[10]), .ZN(n551) );
  INV_X1 U161 ( .A(A[14]), .ZN(n559) );
  INV_X1 U162 ( .A(A[22]), .ZN(n575) );
  INV_X1 U163 ( .A(A[18]), .ZN(n567) );
  NAND2_X1 U164 ( .A1(B[10]), .A2(n551), .ZN(n129) );
  NAND2_X1 U165 ( .A1(B[14]), .A2(n559), .ZN(n117) );
  NAND2_X1 U166 ( .A1(B[22]), .A2(n575), .ZN(n93) );
  NAND2_X1 U167 ( .A1(B[26]), .A2(n583), .ZN(n81) );
  INV_X1 U168 ( .A(A[12]), .ZN(n554) );
  INV_X1 U169 ( .A(A[20]), .ZN(n570) );
  INV_X1 U170 ( .A(A[8]), .ZN(n546) );
  INV_X1 U171 ( .A(A[16]), .ZN(n562) );
  INV_X1 U173 ( .A(A[24]), .ZN(n578) );
  NAND2_X1 U174 ( .A1(B[18]), .A2(n567), .ZN(n105) );
  INV_X1 U175 ( .A(A[4]), .ZN(n538) );
  NAND2_X1 U177 ( .A1(B[7]), .A2(n545), .ZN(n138) );
  INV_X1 U178 ( .A(A[2]), .ZN(n535) );
  NAND2_X1 U179 ( .A1(B[5]), .A2(n540), .ZN(n144) );
  NAND2_X1 U180 ( .A1(B[29]), .A2(n588), .ZN(n72) );
  INV_X1 U181 ( .A(A[6]), .ZN(n543) );
  INV_X1 U182 ( .A(A[0]), .ZN(n533) );
  NAND2_X1 U183 ( .A1(B[6]), .A2(n543), .ZN(n141) );
  INV_X1 U184 ( .A(B[31]), .ZN(n592) );
  AND2_X1 U185 ( .A1(B[4]), .A2(n538), .ZN(n148) );
  INV_X1 U186 ( .A(A[28]), .ZN(n586) );
  AND2_X1 U187 ( .A1(B[8]), .A2(n546), .ZN(n136) );
  AND2_X1 U188 ( .A1(B[16]), .A2(n562), .ZN(n112) );
  AND2_X1 U189 ( .A1(B[24]), .A2(n578), .ZN(n88) );
  AND2_X1 U190 ( .A1(B[12]), .A2(n554), .ZN(n124) );
  AND2_X1 U191 ( .A1(B[20]), .A2(n570), .ZN(n100) );
  AND2_X1 U192 ( .A1(B[28]), .A2(n586), .ZN(n76) );
  INV_X1 U193 ( .A(A[29]), .ZN(n588) );
  INV_X1 U194 ( .A(B[30]), .ZN(n591) );
  OR2_X1 U195 ( .A1(n551), .A2(B[10]), .ZN(n188) );
  OR2_X1 U196 ( .A1(n559), .A2(B[14]), .ZN(n182) );
  OR2_X1 U197 ( .A1(n575), .A2(B[22]), .ZN(n170) );
  OR2_X1 U198 ( .A1(n583), .A2(B[26]), .ZN(n164) );
  OR2_X1 U199 ( .A1(n567), .A2(B[18]), .ZN(n176) );
  OR2_X1 U200 ( .A1(n543), .A2(B[6]), .ZN(n194) );
  OR2_X1 U201 ( .A1(n535), .A2(B[2]), .ZN(n199) );
  INV_X1 U202 ( .A(n202), .ZN(n532) );
  AOI21_X1 U203 ( .B1(A[1]), .B2(n201), .A(n590), .ZN(n202) );
  INV_X1 U204 ( .A(NE), .ZN(EQ) );
  INV_X1 U205 ( .A(GE), .ZN(LT) );
endmodule


module ALU_BEHAVIORAL_NBIT32 ( FUNC, DATA1, DATA2, OUTALU );
  input [3:0] FUNC;
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  wire   N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605,
         N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
  assign N555 = DATA1[0];
  assign N556 = DATA1[1];
  assign N557 = DATA1[2];
  assign N558 = DATA1[3];
  assign N559 = DATA1[4];
  assign N560 = DATA1[5];
  assign N561 = DATA1[6];
  assign N562 = DATA1[7];
  assign N563 = DATA1[8];
  assign N564 = DATA1[9];
  assign N565 = DATA1[10];
  assign N566 = DATA1[11];
  assign N567 = DATA1[12];
  assign N568 = DATA1[13];
  assign N569 = DATA1[14];
  assign N570 = DATA1[15];
  assign N571 = DATA1[16];
  assign N572 = DATA1[17];
  assign N573 = DATA1[18];
  assign N574 = DATA1[19];
  assign N575 = DATA1[20];
  assign N576 = DATA1[21];
  assign N577 = DATA1[22];
  assign N578 = DATA1[23];
  assign N579 = DATA1[24];
  assign N580 = DATA1[25];
  assign N581 = DATA1[26];
  assign N582 = DATA1[27];
  assign N583 = DATA1[28];
  assign N584 = DATA1[29];
  assign N585 = DATA1[30];
  assign N586 = DATA1[31];

  DLH_X1 \OUTALU_reg[31]  ( .G(n1507), .D(N619), .Q(OUTALU[31]) );
  DLH_X1 \OUTALU_reg[30]  ( .G(n1506), .D(N618), .Q(OUTALU[30]) );
  DLH_X1 \OUTALU_reg[29]  ( .G(n1508), .D(N617), .Q(OUTALU[29]) );
  DLH_X1 \OUTALU_reg[28]  ( .G(n1507), .D(N616), .Q(OUTALU[28]) );
  DLH_X1 \OUTALU_reg[27]  ( .G(n1507), .D(N615), .Q(OUTALU[27]) );
  DLH_X1 \OUTALU_reg[26]  ( .G(n1507), .D(N614), .Q(OUTALU[26]) );
  DLH_X1 \OUTALU_reg[25]  ( .G(n1507), .D(N613), .Q(OUTALU[25]) );
  DLH_X1 \OUTALU_reg[24]  ( .G(n1507), .D(N612), .Q(OUTALU[24]) );
  DLH_X1 \OUTALU_reg[23]  ( .G(n1507), .D(N611), .Q(OUTALU[23]) );
  DLH_X1 \OUTALU_reg[22]  ( .G(n1507), .D(N610), .Q(OUTALU[22]) );
  DLH_X1 \OUTALU_reg[21]  ( .G(n1506), .D(N609), .Q(OUTALU[21]) );
  DLH_X1 \OUTALU_reg[20]  ( .G(n1506), .D(N608), .Q(OUTALU[20]) );
  DLH_X1 \OUTALU_reg[19]  ( .G(n1506), .D(N607), .Q(OUTALU[19]) );
  DLH_X1 \OUTALU_reg[18]  ( .G(n1506), .D(N606), .Q(OUTALU[18]) );
  DLH_X1 \OUTALU_reg[17]  ( .G(n1506), .D(N605), .Q(OUTALU[17]) );
  DLH_X1 \OUTALU_reg[16]  ( .G(n1506), .D(N604), .Q(OUTALU[16]) );
  DLH_X1 \OUTALU_reg[15]  ( .G(n1506), .D(N603), .Q(OUTALU[15]) );
  DLH_X1 \OUTALU_reg[14]  ( .G(n1506), .D(N602), .Q(OUTALU[14]) );
  DLH_X1 \OUTALU_reg[13]  ( .G(n1507), .D(N601), .Q(OUTALU[13]) );
  DLH_X1 \OUTALU_reg[12]  ( .G(n1507), .D(N600), .Q(OUTALU[12]) );
  DLH_X1 \OUTALU_reg[11]  ( .G(n1506), .D(N599), .Q(OUTALU[11]) );
  DLH_X1 \OUTALU_reg[10]  ( .G(n1506), .D(N598), .Q(OUTALU[10]) );
  DLH_X1 \OUTALU_reg[9]  ( .G(n1508), .D(N597), .Q(OUTALU[9]) );
  DLH_X1 \OUTALU_reg[8]  ( .G(n1508), .D(N596), .Q(OUTALU[8]) );
  DLH_X1 \OUTALU_reg[7]  ( .G(n1508), .D(N595), .Q(OUTALU[7]) );
  DLH_X1 \OUTALU_reg[6]  ( .G(n1508), .D(N594), .Q(OUTALU[6]) );
  DLH_X1 \OUTALU_reg[5]  ( .G(n1508), .D(N593), .Q(OUTALU[5]) );
  DLH_X1 \OUTALU_reg[4]  ( .G(n1508), .D(N592), .Q(OUTALU[4]) );
  DLH_X1 \OUTALU_reg[3]  ( .G(n1508), .D(N591), .Q(OUTALU[3]) );
  DLH_X1 \OUTALU_reg[2]  ( .G(n1508), .D(N590), .Q(OUTALU[2]) );
  DLH_X1 \OUTALU_reg[1]  ( .G(n1507), .D(N589), .Q(OUTALU[1]) );
  DLH_X1 \OUTALU_reg[0]  ( .G(n1508), .D(N588), .Q(OUTALU[0]) );
  NAND3_X1 U535 ( .A1(n149), .A2(n150), .A3(n1579), .ZN(n148) );
  NAND3_X1 U536 ( .A1(n149), .A2(n174), .A3(n1579), .ZN(n173) );
  NAND3_X1 U537 ( .A1(n317), .A2(n1609), .A3(DATA2[4]), .ZN(n175) );
  NAND3_X1 U538 ( .A1(n320), .A2(n321), .A3(n322), .ZN(N603) );
  NAND3_X1 U539 ( .A1(n441), .A2(n442), .A3(n443), .ZN(N591) );
  NAND3_X1 U540 ( .A1(n456), .A2(n457), .A3(n458), .ZN(N590) );
  OAI33_X1 U541 ( .A1(n369), .A2(n438), .A3(n1572), .B1(n492), .B2(n493), .B3(
        n1612), .ZN(n491) );
  NAND3_X1 U542 ( .A1(n1578), .A2(n1609), .A3(n317), .ZN(n331) );
  NAND3_X1 U543 ( .A1(n317), .A2(FUNC[0]), .A3(DATA2[4]), .ZN(n369) );
  NAND3_X1 U544 ( .A1(FUNC[0]), .A2(n1578), .A3(n317), .ZN(n208) );
  ALU_BEHAVIORAL_NBIT32_DW01_sub_0 sub_31 ( .A({N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555}), .B(DATA2), .CI(1'b0), .DIFF({N452, N451, N450, 
        N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, 
        N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, 
        N425, N424, N423, N422, N421}) );
  ALU_BEHAVIORAL_NBIT32_DW01_add_1 add_30 ( .A({N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555}), .B(DATA2), .CI(1'b0), .SUM({N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389}) );
  ALU_BEHAVIORAL_NBIT32_DW01_cmp6_0 r76 ( .A({N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555}), .B(DATA2), .TC(1'b0), .LT(N551), .GT(N552), .EQ(
        N549), .LE(N553), .GE(N554), .NE(N550) );
  NOR3_X1 U2 ( .A1(n493), .A2(FUNC[0]), .A3(n1612), .ZN(n151) );
  OAI22_X1 U3 ( .A1(n1453), .A2(n1524), .B1(n1454), .B2(n1523), .ZN(n174) );
  NOR2_X1 U4 ( .A1(n369), .A2(n1571), .ZN(n380) );
  NOR2_X2 U8 ( .A1(n1572), .A2(n208), .ZN(n308) );
  OAI221_X1 U9 ( .B1(n1500), .B2(n1523), .C1(n1498), .C2(n1524), .A(n455), 
        .ZN(n209) );
  OAI221_X1 U10 ( .B1(n1501), .B2(n1554), .C1(n1498), .C2(n1552), .A(n480), 
        .ZN(n274) );
  OAI221_X1 U11 ( .B1(n1501), .B2(n1560), .C1(n1498), .C2(n1558), .A(n503), 
        .ZN(n245) );
  OAI221_X1 U12 ( .B1(n1501), .B2(n1562), .C1(n1498), .C2(n1560), .A(n478), 
        .ZN(n233) );
  OAI221_X1 U13 ( .B1(n1500), .B2(n1564), .C1(n1562), .C2(n1495), .A(n464), 
        .ZN(n224) );
  OAI221_X1 U14 ( .B1(n1499), .B2(n1525), .C1(n1497), .C2(n1526), .A(n428), 
        .ZN(n180) );
  OAI221_X1 U15 ( .B1(n1499), .B2(n1526), .C1(n1497), .C2(n1528), .A(n419), 
        .ZN(n158) );
  AND2_X1 U16 ( .A1(DATA2[1]), .A2(n1569), .ZN(n1452) );
  OR2_X1 U17 ( .A1(DATA2[0]), .A2(DATA2[1]), .ZN(n1453) );
  NOR2_X1 U18 ( .A1(n175), .A2(n1571), .ZN(n161) );
  OR2_X1 U19 ( .A1(n1505), .A2(n164), .ZN(n130) );
  INV_X1 U20 ( .A(n1502), .ZN(n1499) );
  INV_X1 U21 ( .A(n1502), .ZN(n1500) );
  INV_X1 U22 ( .A(n1452), .ZN(n1495) );
  INV_X1 U23 ( .A(n1453), .ZN(n1478) );
  INV_X1 U24 ( .A(n1453), .ZN(n1477) );
  INV_X1 U25 ( .A(n1452), .ZN(n1498) );
  INV_X1 U26 ( .A(n1452), .ZN(n1496) );
  INV_X1 U27 ( .A(n1452), .ZN(n1497) );
  INV_X1 U28 ( .A(n149), .ZN(n1572) );
  BUF_X1 U29 ( .A(n123), .Z(n1504) );
  BUF_X1 U30 ( .A(n123), .Z(n1503) );
  BUF_X1 U31 ( .A(n131), .Z(n1489) );
  BUF_X1 U32 ( .A(n131), .Z(n1488) );
  BUF_X1 U33 ( .A(n134), .Z(n1459) );
  BUF_X1 U34 ( .A(n134), .Z(n1460) );
  BUF_X1 U35 ( .A(n123), .Z(n1505) );
  BUF_X1 U36 ( .A(n134), .Z(n1461) );
  BUF_X1 U37 ( .A(n134), .Z(n1462) );
  INV_X1 U38 ( .A(n1491), .ZN(n1490) );
  INV_X1 U39 ( .A(n1481), .ZN(n1480) );
  AOI21_X1 U40 ( .B1(n1479), .B2(n1480), .A(n1491), .ZN(n453) );
  BUF_X1 U41 ( .A(n1608), .Z(n1463) );
  BUF_X1 U42 ( .A(n1608), .Z(n1464) );
  BUF_X1 U43 ( .A(n1466), .Z(n1470) );
  BUF_X1 U44 ( .A(n1465), .Z(n1467) );
  BUF_X1 U45 ( .A(n1465), .Z(n1468) );
  BUF_X1 U46 ( .A(n1465), .Z(n1469) );
  BUF_X1 U47 ( .A(n1466), .Z(n1471) );
  OAI222_X1 U48 ( .A1(n1454), .A2(n1524), .B1(n1495), .B2(n1523), .C1(n1453), 
        .C2(n1525), .ZN(n150) );
  NOR2_X2 U49 ( .A1(n1572), .A2(n331), .ZN(n136) );
  AOI222_X1 U50 ( .A1(n161), .A2(n178), .B1(n1488), .B2(n179), .C1(n157), .C2(
        n180), .ZN(n167) );
  AOI222_X1 U51 ( .A1(n1462), .A2(n155), .B1(n1488), .B2(n156), .C1(n157), 
        .C2(n158), .ZN(n142) );
  AOI222_X1 U52 ( .A1(n1488), .A2(n213), .B1(n1504), .B2(n212), .C1(n1461), 
        .C2(n209), .ZN(n364) );
  AOI222_X1 U53 ( .A1(n1488), .A2(n135), .B1(n1505), .B2(n132), .C1(n157), 
        .C2(n209), .ZN(n202) );
  AOI222_X1 U54 ( .A1(n1579), .A2(n133), .B1(n1462), .B2(n135), .C1(n136), 
        .C2(n137), .ZN(n118) );
  OAI221_X1 U55 ( .B1(n1527), .B2(n242), .C1(n1509), .C2(n1572), .A(n327), 
        .ZN(n133) );
  INV_X1 U56 ( .A(n213), .ZN(n1527) );
  INV_X1 U57 ( .A(n209), .ZN(n1509) );
  AOI22_X1 U58 ( .A1(n328), .A2(n214), .B1(n329), .B2(n212), .ZN(n327) );
  AOI222_X1 U59 ( .A1(n1576), .A2(n299), .B1(n136), .B2(n158), .C1(n1460), 
        .C2(n162), .ZN(n293) );
  AOI222_X1 U60 ( .A1(n1576), .A2(n291), .B1(n136), .B2(n213), .C1(n1462), 
        .C2(n212), .ZN(n285) );
  AOI222_X1 U61 ( .A1(n332), .A2(n255), .B1(n1489), .B2(n209), .C1(n380), .C2(
        n256), .ZN(n404) );
  AOI22_X1 U62 ( .A1(n150), .A2(n1459), .B1(n162), .B2(n1504), .ZN(n378) );
  AOI22_X1 U63 ( .A1(n150), .A2(n136), .B1(n160), .B2(n1504), .ZN(n340) );
  AOI22_X1 U64 ( .A1(n150), .A2(n161), .B1(n155), .B2(n1503), .ZN(n263) );
  AOI22_X1 U65 ( .A1(n150), .A2(n157), .B1(n156), .B2(n1503), .ZN(n221) );
  AOI22_X1 U66 ( .A1(n181), .A2(n1503), .B1(n174), .B2(n136), .ZN(n350) );
  AOI22_X1 U67 ( .A1(n182), .A2(n1503), .B1(n174), .B2(n161), .ZN(n272) );
  AOI22_X1 U68 ( .A1(n209), .A2(n161), .B1(n135), .B2(n1503), .ZN(n252) );
  AOI22_X1 U69 ( .A1(n174), .A2(n1460), .B1(n178), .B2(n1503), .ZN(n389) );
  AOI22_X1 U70 ( .A1(n1460), .A2(n241), .B1(n192), .B2(n1503), .ZN(n399) );
  AOI22_X1 U71 ( .A1(n174), .A2(n159), .B1(n183), .B2(n1503), .ZN(n306) );
  AOI22_X1 U72 ( .A1(n174), .A2(n157), .B1(n179), .B2(n1503), .ZN(n231) );
  NOR2_X1 U73 ( .A1(n1575), .A2(n1573), .ZN(n149) );
  AOI22_X1 U74 ( .A1(n197), .A2(n1503), .B1(n159), .B2(n241), .ZN(n316) );
  AOI22_X1 U75 ( .A1(n194), .A2(n1503), .B1(n157), .B2(n241), .ZN(n240) );
  NAND4_X1 U76 ( .A1(n215), .A2(n216), .A3(n217), .A4(n218), .ZN(N614) );
  AOI222_X1 U77 ( .A1(N415), .A2(n1483), .B1(n1480), .B2(n224), .C1(N447), 
        .C2(n1485), .ZN(n215) );
  AOI222_X1 U78 ( .A1(n1472), .A2(n1565), .B1(n159), .B2(n162), .C1(n136), 
        .C2(n160), .ZN(n216) );
  AOI222_X1 U79 ( .A1(n1461), .A2(n163), .B1(n1488), .B2(n155), .C1(n161), 
        .C2(n158), .ZN(n217) );
  NAND4_X1 U80 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(N613) );
  AOI222_X1 U81 ( .A1(N414), .A2(n1482), .B1(n1480), .B2(n233), .C1(N446), 
        .C2(n1485), .ZN(n225) );
  AOI222_X1 U82 ( .A1(n1472), .A2(n1563), .B1(n159), .B2(n178), .C1(n136), 
        .C2(n181), .ZN(n226) );
  AOI222_X1 U83 ( .A1(n1462), .A2(n183), .B1(n161), .B2(n180), .C1(n1489), 
        .C2(n182), .ZN(n227) );
  NAND4_X1 U84 ( .A1(n234), .A2(n235), .A3(n236), .A4(n237), .ZN(N612) );
  AOI222_X1 U85 ( .A1(N413), .A2(n1483), .B1(n1473), .B2(n1561), .C1(N445), 
        .C2(n1485), .ZN(n234) );
  AOI222_X1 U86 ( .A1(n159), .A2(n192), .B1(n161), .B2(n244), .C1(n1488), .C2(
        n198), .ZN(n236) );
  AOI222_X1 U87 ( .A1(n164), .A2(n245), .B1(n1462), .B2(n197), .C1(n136), .C2(
        n199), .ZN(n235) );
  NAND4_X1 U88 ( .A1(n300), .A2(n301), .A3(n302), .A4(n303), .ZN(N605) );
  AOI222_X1 U89 ( .A1(n1472), .A2(n274), .B1(n308), .B2(n1563), .C1(n1458), 
        .C2(n233), .ZN(n301) );
  AOI222_X1 U90 ( .A1(N406), .A2(n1483), .B1(n1480), .B2(n309), .C1(N438), 
        .C2(n1486), .ZN(n300) );
  AOI222_X1 U91 ( .A1(n1459), .A2(n178), .B1(n136), .B2(n180), .C1(n1489), 
        .C2(n181), .ZN(n302) );
  NAND4_X1 U92 ( .A1(n266), .A2(n267), .A3(n268), .A4(n269), .ZN(N609) );
  AOI222_X1 U93 ( .A1(N410), .A2(n1483), .B1(n1480), .B2(n274), .C1(N442), 
        .C2(n1485), .ZN(n266) );
  AOI222_X1 U94 ( .A1(n1472), .A2(n233), .B1(n1460), .B2(n181), .C1(n1456), 
        .C2(n1563), .ZN(n267) );
  AOI222_X1 U95 ( .A1(n136), .A2(n178), .B1(n1488), .B2(n183), .C1(n159), .C2(
        n180), .ZN(n268) );
  NAND4_X1 U96 ( .A1(n257), .A2(n258), .A3(n259), .A4(n260), .ZN(N610) );
  AOI222_X1 U97 ( .A1(N411), .A2(n1483), .B1(n1473), .B2(n224), .C1(N443), 
        .C2(n1486), .ZN(n257) );
  AOI222_X1 U98 ( .A1(n1457), .A2(n1565), .B1(n136), .B2(n162), .C1(n1480), 
        .C2(n265), .ZN(n258) );
  AOI222_X1 U99 ( .A1(n1460), .A2(n160), .B1(n1488), .B2(n163), .C1(n159), 
        .C2(n158), .ZN(n259) );
  NAND4_X1 U100 ( .A1(n246), .A2(n247), .A3(n248), .A4(n249), .ZN(N611) );
  AOI222_X1 U101 ( .A1(N412), .A2(n1483), .B1(n1473), .B2(n256), .C1(N444), 
        .C2(n1486), .ZN(n246) );
  AOI222_X1 U102 ( .A1(n1455), .A2(n1568), .B1(n136), .B2(n212), .C1(n1480), 
        .C2(n255), .ZN(n247) );
  AOI222_X1 U103 ( .A1(n1459), .A2(n214), .B1(n1488), .B2(n137), .C1(n159), 
        .C2(n213), .ZN(n248) );
  NAND4_X1 U104 ( .A1(n310), .A2(n311), .A3(n312), .A4(n313), .ZN(N604) );
  AOI222_X1 U105 ( .A1(n1472), .A2(n283), .B1(n1480), .B2(n319), .C1(n1455), 
        .C2(n245), .ZN(n311) );
  AOI222_X1 U106 ( .A1(N405), .A2(n1483), .B1(n308), .B2(n1561), .C1(N437), 
        .C2(n1486), .ZN(n310) );
  AOI222_X1 U107 ( .A1(n1461), .A2(n192), .B1(n136), .B2(n244), .C1(n1489), 
        .C2(n199), .ZN(n312) );
  NAND4_X1 U108 ( .A1(n275), .A2(n276), .A3(n277), .A4(n278), .ZN(N608) );
  AOI222_X1 U109 ( .A1(N409), .A2(n1483), .B1(n1473), .B2(n245), .C1(N441), 
        .C2(n1486), .ZN(n275) );
  AOI222_X1 U110 ( .A1(n1458), .A2(n1561), .B1(n1459), .B2(n199), .C1(n1480), 
        .C2(n283), .ZN(n276) );
  AOI222_X1 U111 ( .A1(n136), .A2(n192), .B1(n1505), .B2(n198), .C1(n1489), 
        .C2(n197), .ZN(n277) );
  NAND4_X1 U112 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .ZN(N601) );
  AOI222_X1 U113 ( .A1(n1456), .A2(n274), .B1(n1480), .B2(n352), .C1(n308), 
        .C2(n233), .ZN(n345) );
  AOI222_X1 U114 ( .A1(N402), .A2(n1483), .B1(n1473), .B2(n309), .C1(N434), 
        .C2(n1486), .ZN(n344) );
  AOI222_X1 U115 ( .A1(n332), .A2(n1563), .B1(n1488), .B2(n178), .C1(n1459), 
        .C2(n180), .ZN(n346) );
  NAND4_X1 U116 ( .A1(n334), .A2(n335), .A3(n336), .A4(n337), .ZN(N602) );
  AOI222_X1 U117 ( .A1(n1472), .A2(n342), .B1(n1480), .B2(n343), .C1(n1456), 
        .C2(n265), .ZN(n335) );
  AOI222_X1 U118 ( .A1(N403), .A2(n1483), .B1(n308), .B2(n224), .C1(N435), 
        .C2(n1486), .ZN(n334) );
  AOI222_X1 U119 ( .A1(n332), .A2(n1565), .B1(n1488), .B2(n162), .C1(n1459), 
        .C2(n158), .ZN(n336) );
  NAND4_X1 U120 ( .A1(n353), .A2(n354), .A3(n355), .A4(n356), .ZN(N600) );
  AOI222_X1 U121 ( .A1(n1472), .A2(n319), .B1(n1480), .B2(n361), .C1(n1455), 
        .C2(n283), .ZN(n354) );
  AOI222_X1 U122 ( .A1(N401), .A2(n1483), .B1(n308), .B2(n245), .C1(N433), 
        .C2(n1486), .ZN(n353) );
  AOI222_X1 U123 ( .A1(n332), .A2(n1561), .B1(n1505), .B2(n199), .C1(n1489), 
        .C2(n192), .ZN(n355) );
  NAND4_X1 U124 ( .A1(n412), .A2(n413), .A3(n414), .A4(n415), .ZN(N594) );
  AOI222_X1 U125 ( .A1(n1472), .A2(n382), .B1(n1457), .B2(n343), .C1(n308), 
        .C2(n342), .ZN(n413) );
  AOI222_X1 U126 ( .A1(N395), .A2(n1484), .B1(n1480), .B2(n420), .C1(N427), 
        .C2(n1487), .ZN(n412) );
  AOI222_X1 U127 ( .A1(n332), .A2(n265), .B1(n1489), .B2(n150), .C1(n380), 
        .C2(n224), .ZN(n414) );
  NAND4_X1 U128 ( .A1(n383), .A2(n384), .A3(n385), .A4(n386), .ZN(N597) );
  AOI222_X1 U129 ( .A1(n1457), .A2(n309), .B1(n1473), .B2(n352), .C1(n308), 
        .C2(n274), .ZN(n384) );
  AOI222_X1 U130 ( .A1(N398), .A2(n1484), .B1(n1480), .B2(n392), .C1(N430), 
        .C2(n1486), .ZN(n383) );
  AOI222_X1 U131 ( .A1(n332), .A2(n233), .B1(n1489), .B2(n180), .C1(n380), 
        .C2(n1563), .ZN(n385) );
  NAND4_X1 U132 ( .A1(n372), .A2(n373), .A3(n374), .A4(n375), .ZN(N598) );
  AOI222_X1 U133 ( .A1(n1456), .A2(n342), .B1(n1473), .B2(n343), .C1(n308), 
        .C2(n265), .ZN(n373) );
  AOI222_X1 U134 ( .A1(N399), .A2(n1483), .B1(n1480), .B2(n382), .C1(N431), 
        .C2(n1486), .ZN(n372) );
  AOI222_X1 U135 ( .A1(n332), .A2(n224), .B1(n1488), .B2(n158), .C1(n380), 
        .C2(n1565), .ZN(n374) );
  NAND4_X1 U136 ( .A1(n421), .A2(n422), .A3(n423), .A4(n424), .ZN(N593) );
  AOI222_X1 U137 ( .A1(n1473), .A2(n392), .B1(n1458), .B2(n352), .C1(n308), 
        .C2(n309), .ZN(n422) );
  AOI222_X1 U138 ( .A1(N394), .A2(n1484), .B1(n1480), .B2(n429), .C1(N426), 
        .C2(n1487), .ZN(n421) );
  AOI222_X1 U139 ( .A1(n332), .A2(n274), .B1(n1488), .B2(n174), .C1(n380), 
        .C2(n233), .ZN(n423) );
  NAND4_X1 U140 ( .A1(n393), .A2(n394), .A3(n395), .A4(n396), .ZN(N596) );
  AOI222_X1 U141 ( .A1(n1472), .A2(n361), .B1(n1480), .B2(n401), .C1(n1457), 
        .C2(n319), .ZN(n394) );
  AOI222_X1 U142 ( .A1(N397), .A2(n1484), .B1(n308), .B2(n283), .C1(N429), 
        .C2(n1487), .ZN(n393) );
  AOI222_X1 U143 ( .A1(n332), .A2(n245), .B1(n1489), .B2(n244), .C1(n380), 
        .C2(n1561), .ZN(n395) );
  NOR2_X2 U144 ( .A1(n175), .A2(n1574), .ZN(n159) );
  NOR2_X1 U145 ( .A1(n175), .A2(n242), .ZN(n157) );
  NOR2_X1 U146 ( .A1(n1523), .A2(n1453), .ZN(n241) );
  AOI222_X1 U147 ( .A1(n1457), .A2(n392), .B1(n1505), .B2(n174), .C1(n308), 
        .C2(n352), .ZN(n471) );
  OAI221_X1 U148 ( .B1(n1500), .B2(n1562), .C1(n1497), .C2(n1564), .A(n127), 
        .ZN(n124) );
  NOR2_X1 U149 ( .A1(n1574), .A2(n331), .ZN(n123) );
  NOR2_X1 U150 ( .A1(n1571), .A2(n331), .ZN(n131) );
  NOR2_X1 U151 ( .A1(n242), .A2(n331), .ZN(n134) );
  INV_X1 U152 ( .A(n328), .ZN(n1574) );
  INV_X1 U153 ( .A(n329), .ZN(n1571) );
  INV_X1 U154 ( .A(n175), .ZN(n1579) );
  NOR2_X1 U155 ( .A1(n1453), .A2(n1564), .ZN(n177) );
  NOR2_X1 U156 ( .A1(n1453), .A2(n1566), .ZN(n154) );
  INV_X1 U157 ( .A(n331), .ZN(n1577) );
  INV_X1 U158 ( .A(n408), .ZN(n1568) );
  OAI222_X1 U159 ( .A1(n1547), .A2(n1574), .B1(n1553), .B2(n1571), .C1(n1575), 
        .C2(n207), .ZN(n291) );
  INV_X1 U160 ( .A(n324), .ZN(n1547) );
  INV_X1 U161 ( .A(n255), .ZN(n1553) );
  OAI222_X1 U162 ( .A1(n1495), .A2(n1528), .B1(n1501), .B2(n1530), .C1(n1454), 
        .C2(n1526), .ZN(n468) );
  OAI222_X1 U163 ( .A1(n1495), .A2(n1530), .B1(n1501), .B2(n1531), .C1(n1454), 
        .C2(n1528), .ZN(n452) );
  OAI221_X1 U164 ( .B1(n381), .B2(n1572), .C1(n1559), .C2(n242), .A(n461), 
        .ZN(n299) );
  INV_X1 U165 ( .A(n224), .ZN(n1559) );
  AOI22_X1 U166 ( .A1(n329), .A2(n265), .B1(n328), .B2(n342), .ZN(n461) );
  BUF_X1 U167 ( .A(n223), .Z(n1473) );
  INV_X1 U168 ( .A(n438), .ZN(n1561) );
  BUF_X1 U169 ( .A(n223), .Z(n1472) );
  INV_X1 U170 ( .A(n391), .ZN(n1563) );
  INV_X1 U171 ( .A(n434), .ZN(n1570) );
  INV_X1 U172 ( .A(n381), .ZN(n1565) );
  BUF_X1 U173 ( .A(n254), .Z(n1455) );
  BUF_X1 U174 ( .A(n254), .Z(n1456) );
  INV_X1 U175 ( .A(n152), .ZN(n1608) );
  BUF_X1 U176 ( .A(n254), .Z(n1457) );
  BUF_X1 U177 ( .A(n254), .Z(n1458) );
  BUF_X1 U178 ( .A(n1610), .Z(n1465) );
  INV_X1 U179 ( .A(n459), .ZN(n1532) );
  AOI222_X1 U180 ( .A1(n382), .A2(n1456), .B1(n299), .B2(n1580), .C1(n420), 
        .C2(n1472), .ZN(n459) );
  INV_X1 U181 ( .A(n444), .ZN(n1534) );
  AOI222_X1 U182 ( .A1(n411), .A2(n1472), .B1(n291), .B2(n1580), .C1(n371), 
        .C2(n1455), .ZN(n444) );
  INV_X1 U183 ( .A(n323), .ZN(n1548) );
  AOI222_X1 U184 ( .A1(n324), .A2(n1472), .B1(n255), .B2(n1456), .C1(n256), 
        .C2(n308), .ZN(n323) );
  BUF_X1 U185 ( .A(n1610), .Z(n1466) );
  INV_X1 U186 ( .A(n505), .ZN(n1529) );
  AOI22_X1 U187 ( .A1(n440), .A2(n1472), .B1(n401), .B2(n1455), .ZN(n505) );
  AOI22_X1 U188 ( .A1(N559), .A2(n1474), .B1(N560), .B2(n1478), .ZN(n428) );
  AOI22_X1 U189 ( .A1(N560), .A2(n1474), .B1(N561), .B2(n1478), .ZN(n419) );
  OAI221_X1 U190 ( .B1(n1499), .B2(n1531), .C1(n1497), .C2(n1533), .A(n390), 
        .ZN(n178) );
  AOI22_X1 U191 ( .A1(N563), .A2(n1474), .B1(N564), .B2(n1478), .ZN(n390) );
  OAI221_X1 U192 ( .B1(n1499), .B2(n1530), .C1(n1497), .C2(n1531), .A(n400), 
        .ZN(n192) );
  AOI22_X1 U193 ( .A1(N562), .A2(n1474), .B1(N563), .B2(n1478), .ZN(n400) );
  OAI221_X1 U194 ( .B1(n1499), .B2(n1535), .C1(n1496), .C2(n1536), .A(n370), 
        .ZN(n212) );
  AOI22_X1 U195 ( .A1(N565), .A2(n1474), .B1(N566), .B2(n1478), .ZN(n370) );
  OAI221_X1 U196 ( .B1(n1499), .B2(n1536), .C1(n1496), .C2(n1537), .A(n360), 
        .ZN(n199) );
  AOI22_X1 U197 ( .A1(N566), .A2(n1474), .B1(N567), .B2(n1478), .ZN(n360) );
  OAI221_X1 U198 ( .B1(n1499), .B2(n1538), .C1(n1496), .C2(n1539), .A(n341), 
        .ZN(n160) );
  AOI22_X1 U199 ( .A1(N568), .A2(n1474), .B1(N569), .B2(n1478), .ZN(n341) );
  OAI221_X1 U200 ( .B1(n1500), .B2(n1524), .C1(n1497), .C2(n1525), .A(n437), 
        .ZN(n244) );
  AOI22_X1 U201 ( .A1(N558), .A2(n1474), .B1(N559), .B2(n1478), .ZN(n437) );
  OAI221_X1 U202 ( .B1(n1499), .B2(n1539), .C1(n1496), .C2(n1540), .A(n330), 
        .ZN(n214) );
  AOI22_X1 U203 ( .A1(N569), .A2(n1474), .B1(N570), .B2(n1478), .ZN(n330) );
  OAI221_X1 U204 ( .B1(n125), .B2(n1542), .C1(n1496), .C2(n1543), .A(n298), 
        .ZN(n163) );
  AOI22_X1 U205 ( .A1(N572), .A2(n1475), .B1(N573), .B2(n1477), .ZN(n298) );
  OAI221_X1 U206 ( .B1(n1499), .B2(n1540), .C1(n1496), .C2(n1541), .A(n318), 
        .ZN(n197) );
  AOI22_X1 U207 ( .A1(N570), .A2(n1476), .B1(N571), .B2(n1479), .ZN(n318) );
  OAI221_X1 U208 ( .B1(n1501), .B2(n1541), .C1(n1496), .C2(n1542), .A(n307), 
        .ZN(n183) );
  AOI22_X1 U209 ( .A1(N571), .A2(n1476), .B1(N572), .B2(n1477), .ZN(n307) );
  OAI22_X1 U210 ( .A1(n241), .A2(n1573), .B1(DATA2[2]), .B2(n244), .ZN(n191)
         );
  OAI221_X1 U211 ( .B1(n1500), .B2(n1545), .C1(n1496), .C2(n1546), .A(n273), 
        .ZN(n182) );
  AOI22_X1 U212 ( .A1(N575), .A2(n1476), .B1(N576), .B2(n1477), .ZN(n273) );
  OAI221_X1 U213 ( .B1(n1499), .B2(n1549), .C1(n1495), .C2(n1550), .A(n253), 
        .ZN(n135) );
  AOI22_X1 U214 ( .A1(N577), .A2(n1476), .B1(N578), .B2(n1477), .ZN(n253) );
  OAI221_X1 U215 ( .B1(n1501), .B2(n1546), .C1(n1496), .C2(n1549), .A(n264), 
        .ZN(n155) );
  AOI22_X1 U216 ( .A1(N576), .A2(n1476), .B1(N577), .B2(n1477), .ZN(n264) );
  OAI221_X1 U217 ( .B1(n125), .B2(n1554), .C1(n1495), .C2(n1556), .A(n210), 
        .ZN(n132) );
  AOI22_X1 U218 ( .A1(N581), .A2(n1475), .B1(N582), .B2(n1477), .ZN(n210) );
  OAI221_X1 U219 ( .B1(n125), .B2(n1550), .C1(n1495), .C2(n1551), .A(n243), 
        .ZN(n194) );
  AOI22_X1 U220 ( .A1(N578), .A2(n1475), .B1(N579), .B2(n1477), .ZN(n243) );
  OAI221_X1 U221 ( .B1(n125), .B2(n1551), .C1(n1495), .C2(n1552), .A(n232), 
        .ZN(n179) );
  AOI22_X1 U222 ( .A1(N579), .A2(n1476), .B1(N580), .B2(n1477), .ZN(n232) );
  OAI221_X1 U223 ( .B1(n125), .B2(n1552), .C1(n1495), .C2(n1554), .A(n222), 
        .ZN(n156) );
  AOI22_X1 U224 ( .A1(N580), .A2(n1476), .B1(N581), .B2(n1477), .ZN(n222) );
  AOI221_X1 U225 ( .B1(N567), .B2(n357), .C1(DATA2[12]), .C2(n358), .A(n359), 
        .ZN(n356) );
  OAI21_X1 U226 ( .B1(N567), .B2(n1468), .A(n1463), .ZN(n358) );
  OAI221_X1 U227 ( .B1(DATA2[12]), .B2(n1470), .C1(n1493), .C2(n1588), .A(n129), .ZN(n357) );
  NOR3_X1 U228 ( .A1(n191), .A2(n331), .A3(n1575), .ZN(n359) );
  AOI221_X1 U229 ( .B1(DATA2[8]), .B2(n397), .C1(N563), .C2(n398), .A(n1520), 
        .ZN(n396) );
  OAI21_X1 U230 ( .B1(N563), .B2(n1467), .A(n1463), .ZN(n397) );
  OAI221_X1 U231 ( .B1(DATA2[8]), .B2(n1471), .C1(n1492), .C2(n1584), .A(n129), 
        .ZN(n398) );
  INV_X1 U232 ( .A(n399), .ZN(n1520) );
  AOI221_X1 U233 ( .B1(DATA2[10]), .B2(n376), .C1(N565), .C2(n377), .A(n1511), 
        .ZN(n375) );
  OAI21_X1 U234 ( .B1(N565), .B2(n1468), .A(n1463), .ZN(n376) );
  OAI221_X1 U235 ( .B1(DATA2[10]), .B2(n1471), .C1(n1492), .C2(n1586), .A(n129), .ZN(n377) );
  INV_X1 U236 ( .A(n378), .ZN(n1511) );
  AOI221_X1 U237 ( .B1(DATA2[16]), .B2(n314), .C1(N571), .C2(n315), .A(n1521), 
        .ZN(n313) );
  OAI21_X1 U238 ( .B1(N571), .B2(n1468), .A(n1464), .ZN(n314) );
  OAI221_X1 U239 ( .B1(DATA2[16]), .B2(n1470), .C1(n1493), .C2(n1592), .A(
        n1490), .ZN(n315) );
  INV_X1 U240 ( .A(n316), .ZN(n1521) );
  AOI221_X1 U241 ( .B1(DATA2[21]), .B2(n270), .C1(N576), .C2(n271), .A(n1518), 
        .ZN(n269) );
  OAI21_X1 U242 ( .B1(N576), .B2(n1469), .A(n1464), .ZN(n270) );
  OAI221_X1 U243 ( .B1(DATA2[21]), .B2(n1470), .C1(n1493), .C2(n1597), .A(
        n1490), .ZN(n271) );
  INV_X1 U244 ( .A(n272), .ZN(n1518) );
  AOI221_X1 U245 ( .B1(DATA2[24]), .B2(n238), .C1(N579), .C2(n239), .A(n1522), 
        .ZN(n237) );
  OAI21_X1 U246 ( .B1(N579), .B2(n1468), .A(n1464), .ZN(n238) );
  OAI221_X1 U247 ( .B1(DATA2[24]), .B2(n1470), .C1(n1493), .C2(n1600), .A(
        n1490), .ZN(n239) );
  INV_X1 U248 ( .A(n240), .ZN(n1522) );
  AOI221_X1 U249 ( .B1(DATA2[25]), .B2(n229), .C1(N580), .C2(n230), .A(n1519), 
        .ZN(n228) );
  OAI21_X1 U250 ( .B1(N580), .B2(n1467), .A(n1464), .ZN(n229) );
  OAI221_X1 U251 ( .B1(DATA2[25]), .B2(n1469), .C1(n1494), .C2(n1601), .A(
        n1490), .ZN(n230) );
  INV_X1 U252 ( .A(n231), .ZN(n1519) );
  AOI221_X1 U253 ( .B1(DATA2[26]), .B2(n219), .C1(N581), .C2(n220), .A(n1514), 
        .ZN(n218) );
  OAI21_X1 U254 ( .B1(N581), .B2(n1467), .A(n1464), .ZN(n219) );
  OAI221_X1 U255 ( .B1(DATA2[26]), .B2(n1469), .C1(n1494), .C2(n1602), .A(
        n1490), .ZN(n220) );
  INV_X1 U256 ( .A(n221), .ZN(n1514) );
  AOI221_X1 U257 ( .B1(N560), .B2(n425), .C1(n1504), .C2(n180), .A(n426), .ZN(
        n424) );
  OAI221_X1 U258 ( .B1(DATA2[5]), .B2(n1471), .C1(n1492), .C2(n1581), .A(n129), 
        .ZN(n425) );
  OAI22_X1 U259 ( .A1(n391), .A2(n1570), .B1(n427), .B2(n1581), .ZN(n426) );
  INV_X1 U260 ( .A(DATA2[5]), .ZN(n1581) );
  AOI221_X1 U261 ( .B1(N561), .B2(n416), .C1(n1504), .C2(n158), .A(n417), .ZN(
        n415) );
  OAI221_X1 U262 ( .B1(DATA2[6]), .B2(n1471), .C1(n1492), .C2(n1582), .A(n129), 
        .ZN(n416) );
  OAI22_X1 U263 ( .A1(n381), .A2(n1570), .B1(n418), .B2(n1582), .ZN(n417) );
  INV_X1 U264 ( .A(DATA2[6]), .ZN(n1582) );
  AOI22_X1 U265 ( .A1(n332), .A2(n1568), .B1(n1480), .B2(n333), .ZN(n320) );
  AOI221_X1 U266 ( .B1(N436), .B2(n1487), .C1(N404), .C2(n1482), .A(n1548), 
        .ZN(n322) );
  AOI222_X1 U267 ( .A1(n1577), .A2(n133), .B1(DATA2[15]), .B2(n325), .C1(N570), 
        .C2(n326), .ZN(n321) );
  AOI221_X1 U268 ( .B1(n434), .B2(n1561), .C1(DATA2[4]), .C2(n435), .A(n436), 
        .ZN(n433) );
  OAI21_X1 U269 ( .B1(N559), .B2(n1467), .A(n1463), .ZN(n435) );
  NOR3_X1 U270 ( .A1(n191), .A2(DATA2[3]), .A3(n331), .ZN(n436) );
  AOI221_X1 U271 ( .B1(N575), .B2(n279), .C1(DATA2[20]), .C2(n280), .A(n281), 
        .ZN(n278) );
  OAI21_X1 U272 ( .B1(N575), .B2(n1468), .A(n1464), .ZN(n280) );
  OAI221_X1 U273 ( .B1(DATA2[20]), .B2(n1470), .C1(n1493), .C2(n1596), .A(
        n1490), .ZN(n279) );
  NOR3_X1 U274 ( .A1(n191), .A2(DATA2[3]), .A3(n175), .ZN(n281) );
  AOI221_X1 U275 ( .B1(n1504), .B2(n188), .C1(DATA2[28]), .C2(n189), .A(n190), 
        .ZN(n187) );
  OAI21_X1 U276 ( .B1(N583), .B2(n1467), .A(n1608), .ZN(n189) );
  OAI222_X1 U277 ( .A1(n1495), .A2(n1558), .B1(n1501), .B2(n1556), .C1(n1454), 
        .C2(n1560), .ZN(n188) );
  NOR3_X1 U278 ( .A1(n191), .A2(n1575), .A3(n175), .ZN(n190) );
  AOI22_X1 U279 ( .A1(N557), .A2(n1476), .B1(N558), .B2(n1477), .ZN(n455) );
  OAI221_X1 U280 ( .B1(n1499), .B2(n1528), .C1(n1497), .C2(n1530), .A(n410), 
        .ZN(n213) );
  AOI22_X1 U281 ( .A1(N561), .A2(n1474), .B1(N562), .B2(n1478), .ZN(n410) );
  OAI221_X1 U282 ( .B1(n125), .B2(n1544), .C1(n1496), .C2(n1545), .A(n282), 
        .ZN(n198) );
  AOI22_X1 U283 ( .A1(N574), .A2(n1476), .B1(N575), .B2(n1477), .ZN(n282) );
  OAI221_X1 U284 ( .B1(n1499), .B2(n1537), .C1(n1496), .C2(n1538), .A(n351), 
        .ZN(n181) );
  AOI22_X1 U285 ( .A1(N567), .A2(n1474), .B1(N568), .B2(n1478), .ZN(n351) );
  OAI221_X1 U286 ( .B1(n1499), .B2(n1533), .C1(n1496), .C2(n1535), .A(n379), 
        .ZN(n162) );
  AOI22_X1 U287 ( .A1(N564), .A2(n1474), .B1(N565), .B2(n1478), .ZN(n379) );
  OAI221_X1 U288 ( .B1(n125), .B2(n1543), .C1(n1496), .C2(n1544), .A(n290), 
        .ZN(n137) );
  AOI22_X1 U289 ( .A1(N573), .A2(n1476), .B1(N574), .B2(n1477), .ZN(n290) );
  INV_X1 U290 ( .A(DATA2[3]), .ZN(n1575) );
  INV_X1 U291 ( .A(DATA2[0]), .ZN(n1569) );
  NAND2_X1 U292 ( .A1(DATA2[1]), .A2(DATA2[0]), .ZN(n125) );
  NAND4_X1 U293 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(N615) );
  AOI221_X1 U294 ( .B1(N582), .B2(n204), .C1(DATA2[27]), .C2(n205), .A(n206), 
        .ZN(n203) );
  AOI222_X1 U295 ( .A1(N416), .A2(n1482), .B1(n136), .B2(n214), .C1(N448), 
        .C2(n1485), .ZN(n200) );
  AOI222_X1 U296 ( .A1(n159), .A2(n212), .B1(n161), .B2(n213), .C1(n1460), 
        .C2(n137), .ZN(n201) );
  NAND4_X1 U297 ( .A1(n140), .A2(n141), .A3(n142), .A4(n143), .ZN(N618) );
  AOI222_X1 U298 ( .A1(N419), .A2(n1482), .B1(n1480), .B2(n1565), .C1(N451), 
        .C2(n1485), .ZN(n140) );
  AOI221_X1 U299 ( .B1(N585), .B2(n144), .C1(n1504), .C2(n145), .A(n146), .ZN(
        n143) );
  AOI222_X1 U300 ( .A1(n159), .A2(n160), .B1(n161), .B2(n162), .C1(n136), .C2(
        n163), .ZN(n141) );
  NAND4_X1 U301 ( .A1(n184), .A2(n185), .A3(n186), .A4(n187), .ZN(N616) );
  AOI222_X1 U302 ( .A1(N417), .A2(n1482), .B1(n1480), .B2(n1561), .C1(N449), 
        .C2(n1485), .ZN(n184) );
  AOI222_X1 U303 ( .A1(n161), .A2(n192), .B1(N583), .B2(n193), .C1(n1489), 
        .C2(n194), .ZN(n186) );
  AOI222_X1 U304 ( .A1(n136), .A2(n197), .B1(n1461), .B2(n198), .C1(n159), 
        .C2(n199), .ZN(n185) );
  NAND4_X1 U305 ( .A1(n165), .A2(n166), .A3(n167), .A4(n168), .ZN(N617) );
  AOI222_X1 U306 ( .A1(N418), .A2(n1482), .B1(n1480), .B2(n1563), .C1(N450), 
        .C2(n1485), .ZN(n165) );
  AOI221_X1 U307 ( .B1(N584), .B2(n169), .C1(n1504), .C2(n170), .A(n171), .ZN(
        n168) );
  AOI222_X1 U308 ( .A1(n159), .A2(n181), .B1(n1461), .B2(n182), .C1(n136), 
        .C2(n183), .ZN(n166) );
  NAND4_X1 U309 ( .A1(n117), .A2(n118), .A3(n119), .A4(n120), .ZN(N619) );
  AOI22_X1 U310 ( .A1(N452), .A2(n1485), .B1(N420), .B2(n1482), .ZN(n117) );
  AOI222_X1 U311 ( .A1(N586), .A2(n121), .B1(DATA2[31]), .B2(n122), .C1(n1505), 
        .C2(n124), .ZN(n120) );
  AOI22_X1 U312 ( .A1(n1568), .A2(n130), .B1(n1489), .B2(n132), .ZN(n119) );
  NAND4_X1 U313 ( .A1(n292), .A2(n293), .A3(n294), .A4(n295), .ZN(N606) );
  AOI22_X1 U314 ( .A1(N439), .A2(n1485), .B1(N407), .B2(n1482), .ZN(n292) );
  AOI22_X1 U315 ( .A1(n159), .A2(n150), .B1(n1489), .B2(n160), .ZN(n294) );
  AOI222_X1 U316 ( .A1(n1504), .A2(n163), .B1(DATA2[18]), .B2(n296), .C1(N573), 
        .C2(n297), .ZN(n295) );
  NAND4_X1 U317 ( .A1(n284), .A2(n285), .A3(n286), .A4(n287), .ZN(N607) );
  AOI22_X1 U318 ( .A1(N440), .A2(n1485), .B1(N408), .B2(n1482), .ZN(n284) );
  AOI222_X1 U319 ( .A1(n1504), .A2(n137), .B1(DATA2[19]), .B2(n288), .C1(N574), 
        .C2(n289), .ZN(n287) );
  AOI22_X1 U320 ( .A1(n159), .A2(n209), .B1(n1489), .B2(n214), .ZN(n286) );
  NAND4_X1 U321 ( .A1(n362), .A2(n363), .A3(n364), .A4(n365), .ZN(N599) );
  AOI222_X1 U322 ( .A1(n1458), .A2(n324), .B1(n1473), .B2(n333), .C1(n308), 
        .C2(n255), .ZN(n363) );
  AOI222_X1 U323 ( .A1(N400), .A2(n1483), .B1(n1480), .B2(n371), .C1(N432), 
        .C2(n1486), .ZN(n362) );
  AOI221_X1 U324 ( .B1(N566), .B2(n366), .C1(DATA2[11]), .C2(n367), .A(n368), 
        .ZN(n365) );
  NAND4_X1 U325 ( .A1(n402), .A2(n403), .A3(n404), .A4(n405), .ZN(N595) );
  AOI222_X1 U326 ( .A1(n1480), .A2(n411), .B1(n1458), .B2(n333), .C1(n308), 
        .C2(n324), .ZN(n403) );
  AOI222_X1 U327 ( .A1(N396), .A2(n1484), .B1(n1473), .B2(n371), .C1(N428), 
        .C2(n1486), .ZN(n402) );
  AOI221_X1 U328 ( .B1(N562), .B2(n406), .C1(n1504), .C2(n213), .A(n407), .ZN(
        n405) );
  OR2_X1 U329 ( .A1(n1569), .A2(DATA2[1]), .ZN(n1454) );
  OAI21_X1 U330 ( .B1(n147), .B2(n1606), .A(n148), .ZN(n146) );
  AOI21_X1 U331 ( .B1(n151), .B2(n1566), .A(n152), .ZN(n147) );
  NAND4_X1 U332 ( .A1(n430), .A2(n431), .A3(n432), .A4(n433), .ZN(N592) );
  AOI222_X1 U333 ( .A1(n1455), .A2(n361), .B1(n1480), .B2(n440), .C1(n1473), 
        .C2(n401), .ZN(n431) );
  AOI222_X1 U334 ( .A1(n332), .A2(n283), .B1(N559), .B2(n439), .C1(n380), .C2(
        n245), .ZN(n432) );
  AOI222_X1 U335 ( .A1(N393), .A2(n1484), .B1(n308), .B2(n319), .C1(N425), 
        .C2(n1487), .ZN(n430) );
  AOI221_X1 U336 ( .B1(DATA2[14]), .B2(n338), .C1(N569), .C2(n339), .A(n1512), 
        .ZN(n337) );
  OAI21_X1 U337 ( .B1(N569), .B2(n1468), .A(n1463), .ZN(n338) );
  OAI221_X1 U338 ( .B1(DATA2[14]), .B2(n1470), .C1(n1493), .C2(n1590), .A(n129), .ZN(n339) );
  INV_X1 U339 ( .A(n340), .ZN(n1512) );
  AOI221_X1 U340 ( .B1(DATA2[22]), .B2(n261), .C1(N577), .C2(n262), .A(n1513), 
        .ZN(n260) );
  OAI21_X1 U341 ( .B1(N577), .B2(n1468), .A(n1464), .ZN(n261) );
  OAI221_X1 U342 ( .B1(DATA2[22]), .B2(n1469), .C1(n1493), .C2(n1598), .A(
        n1490), .ZN(n262) );
  INV_X1 U343 ( .A(n263), .ZN(n1513) );
  AOI221_X1 U344 ( .B1(DATA2[13]), .B2(n348), .C1(N568), .C2(n349), .A(n1516), 
        .ZN(n347) );
  OAI21_X1 U345 ( .B1(N568), .B2(n1467), .A(n1463), .ZN(n348) );
  OAI221_X1 U346 ( .B1(DATA2[13]), .B2(n1470), .C1(n1493), .C2(n1589), .A(n129), .ZN(n349) );
  INV_X1 U347 ( .A(n350), .ZN(n1516) );
  AOI221_X1 U348 ( .B1(N424), .B2(n1487), .C1(N392), .C2(n1482), .A(n1534), 
        .ZN(n443) );
  AOI222_X1 U349 ( .A1(DATA2[3]), .A2(n450), .B1(N558), .B2(n451), .C1(n1480), 
        .C2(n452), .ZN(n442) );
  AOI22_X1 U350 ( .A1(n1504), .A2(n209), .B1(n308), .B2(n333), .ZN(n441) );
  AOI221_X1 U351 ( .B1(DATA2[23]), .B2(n250), .C1(N578), .C2(n251), .A(n1510), 
        .ZN(n249) );
  OAI21_X1 U352 ( .B1(N578), .B2(n1468), .A(n1464), .ZN(n250) );
  OAI221_X1 U353 ( .B1(DATA2[23]), .B2(n1470), .C1(n1493), .C2(n1599), .A(
        n1490), .ZN(n251) );
  INV_X1 U354 ( .A(n252), .ZN(n1510) );
  AOI221_X1 U355 ( .B1(DATA2[9]), .B2(n387), .C1(N564), .C2(n388), .A(n1515), 
        .ZN(n386) );
  OAI21_X1 U356 ( .B1(N564), .B2(n1467), .A(n1463), .ZN(n387) );
  OAI221_X1 U357 ( .B1(DATA2[9]), .B2(n1471), .C1(n1492), .C2(n1585), .A(n1490), .ZN(n388) );
  INV_X1 U358 ( .A(n389), .ZN(n1515) );
  AOI221_X1 U359 ( .B1(DATA2[17]), .B2(n304), .C1(N572), .C2(n305), .A(n1517), 
        .ZN(n303) );
  OAI21_X1 U360 ( .B1(N572), .B2(n1468), .A(n1464), .ZN(n304) );
  OAI221_X1 U361 ( .B1(DATA2[17]), .B2(n1470), .C1(n1493), .C2(n1593), .A(
        n1490), .ZN(n305) );
  INV_X1 U362 ( .A(n306), .ZN(n1517) );
  AOI221_X1 U363 ( .B1(N555), .B2(n500), .C1(n241), .C2(n130), .A(n501), .ZN(
        n487) );
  OAI221_X1 U364 ( .B1(DATA2[0]), .B2(n1469), .C1(n1492), .C2(n1569), .A(n1490), .ZN(n500) );
  OAI22_X1 U365 ( .A1(n502), .A2(n1481), .B1(n1555), .B2(n1570), .ZN(n501) );
  INV_X1 U366 ( .A(n245), .ZN(n1555) );
  OAI221_X1 U367 ( .B1(n1495), .B2(n1560), .C1(n1454), .C2(n1562), .A(n176), 
        .ZN(n170) );
  AOI21_X1 U368 ( .B1(N581), .B2(n1502), .A(n177), .ZN(n176) );
  OAI221_X1 U369 ( .B1(n1562), .B2(n1495), .C1(n1454), .C2(n1564), .A(n153), 
        .ZN(n145) );
  AOI21_X1 U370 ( .B1(N582), .B2(n1502), .A(n154), .ZN(n153) );
  NOR2_X1 U371 ( .A1(DATA2[2]), .A2(DATA2[3]), .ZN(n328) );
  NOR2_X1 U372 ( .A1(n1573), .A2(DATA2[3]), .ZN(n329) );
  NAND2_X1 U373 ( .A1(DATA2[3]), .A2(n1573), .ZN(n242) );
  INV_X1 U374 ( .A(N584), .ZN(n1564) );
  INV_X1 U375 ( .A(N583), .ZN(n1562) );
  INV_X1 U376 ( .A(DATA2[2]), .ZN(n1573) );
  INV_X1 U377 ( .A(N556), .ZN(n1524) );
  INV_X1 U378 ( .A(N562), .ZN(n1533) );
  INV_X1 U379 ( .A(N561), .ZN(n1531) );
  INV_X1 U380 ( .A(N560), .ZN(n1530) );
  AOI221_X1 U381 ( .B1(N423), .B2(n1487), .C1(N391), .C2(n1482), .A(n1532), 
        .ZN(n458) );
  AOI222_X1 U382 ( .A1(DATA2[2]), .A2(n466), .B1(N557), .B2(n467), .C1(n1480), 
        .C2(n468), .ZN(n457) );
  AOI22_X1 U383 ( .A1(n1504), .A2(n150), .B1(n308), .B2(n343), .ZN(n456) );
  INV_X1 U384 ( .A(N575), .ZN(n1549) );
  INV_X1 U385 ( .A(N567), .ZN(n1539) );
  INV_X1 U386 ( .A(N566), .ZN(n1538) );
  INV_X1 U387 ( .A(N578), .ZN(n1552) );
  INV_X1 U388 ( .A(N568), .ZN(n1540) );
  INV_X1 U389 ( .A(N564), .ZN(n1536) );
  INV_X1 U390 ( .A(N576), .ZN(n1550) );
  INV_X1 U391 ( .A(N577), .ZN(n1551) );
  INV_X1 U392 ( .A(N565), .ZN(n1537) );
  INV_X1 U393 ( .A(N569), .ZN(n1541) );
  INV_X1 U394 ( .A(N563), .ZN(n1535) );
  INV_X1 U395 ( .A(N571), .ZN(n1543) );
  INV_X1 U396 ( .A(N572), .ZN(n1544) );
  INV_X1 U397 ( .A(N579), .ZN(n1554) );
  INV_X1 U398 ( .A(N558), .ZN(n1526) );
  INV_X1 U399 ( .A(N574), .ZN(n1546) );
  INV_X1 U400 ( .A(N573), .ZN(n1545) );
  INV_X1 U401 ( .A(N570), .ZN(n1542) );
  INV_X1 U402 ( .A(N580), .ZN(n1556) );
  INV_X1 U403 ( .A(N582), .ZN(n1560) );
  INV_X1 U404 ( .A(N559), .ZN(n1528) );
  INV_X1 U405 ( .A(N557), .ZN(n1525) );
  INV_X1 U406 ( .A(N555), .ZN(n1523) );
  INV_X1 U407 ( .A(N581), .ZN(n1558) );
  INV_X1 U408 ( .A(N585), .ZN(n1566) );
  NAND2_X1 U409 ( .A1(n1479), .A2(N586), .ZN(n408) );
  NAND2_X1 U410 ( .A1(N585), .A2(n1476), .ZN(n127) );
  NAND4_X1 U411 ( .A1(n470), .A2(n471), .A3(n472), .A4(n473), .ZN(N589) );
  AOI211_X1 U412 ( .C1(N556), .C2(n474), .A(n475), .B(n476), .ZN(n473) );
  AOI222_X1 U413 ( .A1(n332), .A2(n309), .B1(DATA2[1]), .B2(n479), .C1(n380), 
        .C2(n274), .ZN(n472) );
  AOI222_X1 U414 ( .A1(N390), .A2(n1484), .B1(n1473), .B2(n429), .C1(N422), 
        .C2(n1487), .ZN(n470) );
  OAI221_X1 U415 ( .B1(DATA2[28]), .B2(n1469), .C1(n1494), .C2(n1604), .A(n195), .ZN(n193) );
  INV_X1 U416 ( .A(DATA2[28]), .ZN(n1604) );
  AOI21_X1 U417 ( .B1(n1479), .B2(n1503), .A(n1491), .ZN(n195) );
  INV_X1 U418 ( .A(DATA2[4]), .ZN(n1578) );
  OAI21_X1 U419 ( .B1(n172), .B2(n1605), .A(n173), .ZN(n171) );
  AOI21_X1 U420 ( .B1(n151), .B2(n1564), .A(n152), .ZN(n172) );
  AOI22_X1 U421 ( .A1(N580), .A2(n1475), .B1(N579), .B2(n1479), .ZN(n503) );
  AOI22_X1 U422 ( .A1(N581), .A2(n1475), .B1(N580), .B2(n1479), .ZN(n478) );
  AOI22_X1 U423 ( .A1(N582), .A2(n1475), .B1(N581), .B2(n1479), .ZN(n464) );
  AOI22_X1 U424 ( .A1(N577), .A2(n1475), .B1(N576), .B2(n1479), .ZN(n480) );
  OAI221_X1 U425 ( .B1(n1501), .B2(n1552), .C1(n1498), .C2(n1551), .A(n509), 
        .ZN(n283) );
  AOI22_X1 U426 ( .A1(N576), .A2(n1475), .B1(N575), .B2(n1479), .ZN(n509) );
  OAI221_X1 U427 ( .B1(n1501), .B2(n1546), .C1(n1498), .C2(n1545), .A(n508), 
        .ZN(n319) );
  AOI22_X1 U428 ( .A1(N572), .A2(n1476), .B1(N571), .B2(n1479), .ZN(n508) );
  OAI221_X1 U429 ( .B1(n1500), .B2(n1556), .C1(n1498), .C2(n1554), .A(n463), 
        .ZN(n265) );
  AOI22_X1 U430 ( .A1(N578), .A2(n1475), .B1(N577), .B2(n1479), .ZN(n463) );
  OAI221_X1 U431 ( .B1(n1501), .B2(n1549), .C1(n1498), .C2(n1546), .A(n481), 
        .ZN(n309) );
  AOI22_X1 U432 ( .A1(N573), .A2(n1475), .B1(N572), .B2(n1479), .ZN(n481) );
  OAI221_X1 U433 ( .B1(n1500), .B2(n1558), .C1(n1497), .C2(n1556), .A(n447), 
        .ZN(n255) );
  AOI22_X1 U434 ( .A1(N579), .A2(n1475), .B1(N578), .B2(n1479), .ZN(n447) );
  NOR2_X1 U435 ( .A1(n1609), .A2(n1492), .ZN(n152) );
  NOR2_X2 U436 ( .A1(n369), .A2(n1574), .ZN(n332) );
  OAI221_X1 U437 ( .B1(n1500), .B2(n1545), .C1(n1497), .C2(n1544), .A(n454), 
        .ZN(n333) );
  AOI22_X1 U438 ( .A1(N571), .A2(n1475), .B1(N570), .B2(n1477), .ZN(n454) );
  OAI221_X1 U439 ( .B1(n1501), .B2(n1544), .C1(n1498), .C2(n1543), .A(n469), 
        .ZN(n343) );
  AOI22_X1 U440 ( .A1(N570), .A2(n1475), .B1(N569), .B2(n1479), .ZN(n469) );
  OAI221_X1 U441 ( .B1(n1501), .B2(n1543), .C1(n1498), .C2(n1542), .A(n482), 
        .ZN(n352) );
  AOI22_X1 U442 ( .A1(N569), .A2(n1475), .B1(N568), .B2(n1479), .ZN(n482) );
  AOI211_X1 U443 ( .C1(n1452), .C2(N586), .A(n1567), .B(n177), .ZN(n391) );
  INV_X1 U444 ( .A(n127), .ZN(n1567) );
  OAI221_X1 U445 ( .B1(n125), .B2(n1542), .C1(n1495), .C2(n1541), .A(n510), 
        .ZN(n361) );
  AOI22_X1 U446 ( .A1(N568), .A2(n1476), .B1(N567), .B2(n1477), .ZN(n510) );
  OAI221_X1 U447 ( .B1(n1500), .B2(n1550), .C1(n1498), .C2(n1549), .A(n462), 
        .ZN(n342) );
  AOI22_X1 U448 ( .A1(N574), .A2(n1475), .B1(N573), .B2(n1479), .ZN(n462) );
  OAI221_X1 U449 ( .B1(n1566), .B2(n1501), .C1(n1497), .C2(n1564), .A(n446), 
        .ZN(n256) );
  AOI22_X1 U450 ( .A1(N583), .A2(n1475), .B1(N582), .B2(n1479), .ZN(n446) );
  OAI221_X1 U451 ( .B1(n1500), .B2(n1551), .C1(n1497), .C2(n1550), .A(n448), 
        .ZN(n324) );
  AOI22_X1 U452 ( .A1(N575), .A2(n1475), .B1(N574), .B2(n1477), .ZN(n448) );
  OAI221_X1 U453 ( .B1(n1501), .B2(n1539), .C1(n1498), .C2(n1538), .A(n483), 
        .ZN(n392) );
  AOI22_X1 U454 ( .A1(N565), .A2(n1475), .B1(N564), .B2(n1479), .ZN(n483) );
  OAI221_X1 U455 ( .B1(n1501), .B2(n1540), .C1(n1498), .C2(n1539), .A(n465), 
        .ZN(n382) );
  AOI22_X1 U456 ( .A1(N566), .A2(n1475), .B1(N565), .B2(n1479), .ZN(n465) );
  OAI221_X1 U457 ( .B1(n1500), .B2(n1541), .C1(n1497), .C2(n1540), .A(n445), 
        .ZN(n371) );
  AOI22_X1 U458 ( .A1(N567), .A2(n1475), .B1(N566), .B2(n1479), .ZN(n445) );
  OAI221_X1 U459 ( .B1(n1501), .B2(n1538), .C1(n1498), .C2(n1537), .A(n506), 
        .ZN(n401) );
  AOI22_X1 U460 ( .A1(N564), .A2(n1475), .B1(N563), .B2(n1479), .ZN(n506) );
  AOI221_X1 U461 ( .B1(n1502), .B2(N586), .C1(N585), .C2(n1452), .A(n494), 
        .ZN(n438) );
  OAI22_X1 U462 ( .A1(n1564), .A2(n1454), .B1(n1453), .B2(n1562), .ZN(n494) );
  OAI22_X1 U463 ( .A1(DATA2[2]), .A2(n256), .B1(n1568), .B2(n1573), .ZN(n207)
         );
  AOI222_X1 U464 ( .A1(N556), .A2(n1476), .B1(N558), .B2(n1502), .C1(N557), 
        .C2(n1452), .ZN(n502) );
  OAI221_X1 U465 ( .B1(n1501), .B2(n1535), .C1(n1498), .C2(n1533), .A(n484), 
        .ZN(n429) );
  AOI22_X1 U466 ( .A1(N561), .A2(n1475), .B1(N560), .B2(n1479), .ZN(n484) );
  OAI221_X1 U467 ( .B1(n1501), .B2(n1533), .C1(n1496), .C2(n1531), .A(n507), 
        .ZN(n440) );
  AOI22_X1 U468 ( .A1(N560), .A2(n1475), .B1(N559), .B2(n1479), .ZN(n507) );
  OAI221_X1 U469 ( .B1(n1500), .B2(n1537), .C1(n1497), .C2(n1536), .A(n449), 
        .ZN(n411) );
  AOI22_X1 U470 ( .A1(N563), .A2(n1475), .B1(N562), .B2(n1477), .ZN(n449) );
  OAI221_X1 U471 ( .B1(n1500), .B2(n1536), .C1(n1498), .C2(n1535), .A(n460), 
        .ZN(n420) );
  AOI22_X1 U472 ( .A1(N562), .A2(n1475), .B1(N561), .B2(n1479), .ZN(n460) );
  AOI21_X1 U473 ( .B1(n1476), .B2(N586), .A(n154), .ZN(n381) );
  NOR3_X1 U474 ( .A1(n369), .A2(DATA2[3]), .A3(n207), .ZN(n368) );
  NOR3_X1 U475 ( .A1(n369), .A2(n391), .A3(n1572), .ZN(n476) );
  NOR2_X1 U476 ( .A1(n369), .A2(n242), .ZN(n434) );
  NOR3_X1 U477 ( .A1(n207), .A2(DATA2[3]), .A3(n208), .ZN(n206) );
  OAI22_X1 U478 ( .A1(n408), .A2(n1570), .B1(n409), .B2(n1583), .ZN(n407) );
  AOI21_X1 U479 ( .B1(n151), .B2(n1533), .A(n152), .ZN(n409) );
  OAI221_X1 U480 ( .B1(N556), .B2(n1471), .C1(n1492), .C2(n1524), .A(n1463), 
        .ZN(n479) );
  OAI221_X1 U481 ( .B1(DATA2[4]), .B2(n1471), .C1(n1492), .C2(n1578), .A(n1490), .ZN(n439) );
  OAI221_X1 U482 ( .B1(DATA2[15]), .B2(n1470), .C1(n1493), .C2(n1591), .A(
        n1490), .ZN(n326) );
  INV_X1 U483 ( .A(DATA2[15]), .ZN(n1591) );
  OAI221_X1 U484 ( .B1(DATA2[18]), .B2(n1470), .C1(n1493), .C2(n1594), .A(
        n1490), .ZN(n297) );
  INV_X1 U485 ( .A(DATA2[18]), .ZN(n1594) );
  OAI221_X1 U486 ( .B1(DATA2[19]), .B2(n1470), .C1(n1493), .C2(n1595), .A(
        n1490), .ZN(n289) );
  INV_X1 U487 ( .A(DATA2[19]), .ZN(n1595) );
  OAI221_X1 U488 ( .B1(N557), .B2(n1471), .C1(n1492), .C2(n1525), .A(n1463), 
        .ZN(n466) );
  OAI221_X1 U489 ( .B1(N558), .B2(n1471), .C1(n1492), .C2(n1526), .A(n1463), 
        .ZN(n450) );
  OAI221_X1 U490 ( .B1(DATA2[31]), .B2(n1469), .C1(n1494), .C2(n1607), .A(n129), .ZN(n121) );
  INV_X1 U491 ( .A(DATA2[31]), .ZN(n1607) );
  BUF_X1 U492 ( .A(n139), .Z(n1483) );
  OAI221_X1 U493 ( .B1(DATA2[7]), .B2(n1471), .C1(n1492), .C2(n1583), .A(n1490), .ZN(n406) );
  OAI221_X1 U494 ( .B1(DATA2[11]), .B2(n1470), .C1(n1492), .C2(n1587), .A(
        n1490), .ZN(n366) );
  INV_X1 U495 ( .A(DATA2[11]), .ZN(n1587) );
  OAI221_X1 U496 ( .B1(DATA2[27]), .B2(n1469), .C1(n1494), .C2(n1603), .A(n129), .ZN(n204) );
  INV_X1 U497 ( .A(DATA2[27]), .ZN(n1603) );
  OAI221_X1 U498 ( .B1(DATA2[29]), .B2(n1469), .C1(n1494), .C2(n1605), .A(n129), .ZN(n169) );
  OAI221_X1 U499 ( .B1(DATA2[30]), .B2(n1469), .C1(n1494), .C2(n1606), .A(n129), .ZN(n144) );
  NOR2_X1 U500 ( .A1(n242), .A2(n208), .ZN(n254) );
  OAI22_X1 U501 ( .A1(n477), .A2(n1481), .B1(n1557), .B2(n1570), .ZN(n475) );
  INV_X1 U502 ( .A(n233), .ZN(n1557) );
  AOI222_X1 U503 ( .A1(N557), .A2(n1476), .B1(N559), .B2(n1502), .C1(N558), 
        .C2(n1452), .ZN(n477) );
  BUF_X1 U504 ( .A(n138), .Z(n1485) );
  BUF_X1 U505 ( .A(n139), .Z(n1482) );
  BUF_X1 U506 ( .A(n128), .Z(n1492) );
  BUF_X1 U507 ( .A(n138), .Z(n1486) );
  BUF_X1 U508 ( .A(n128), .Z(n1493) );
  NOR2_X1 U509 ( .A1(n208), .A2(n1574), .ZN(n164) );
  NOR2_X1 U510 ( .A1(n1571), .A2(n208), .ZN(n223) );
  BUF_X1 U511 ( .A(n138), .Z(n1487) );
  OAI21_X1 U512 ( .B1(DATA2[3]), .B2(n1467), .A(n453), .ZN(n451) );
  INV_X1 U513 ( .A(n369), .ZN(n1580) );
  BUF_X1 U514 ( .A(n139), .Z(n1484) );
  AOI21_X1 U515 ( .B1(n151), .B2(n1530), .A(n152), .ZN(n427) );
  AOI21_X1 U516 ( .B1(n151), .B2(n1531), .A(n152), .ZN(n418) );
  AOI21_X1 U517 ( .B1(n1609), .B2(n504), .A(n152), .ZN(n129) );
  INV_X1 U518 ( .A(n208), .ZN(n1576) );
  OAI21_X1 U519 ( .B1(N586), .B2(n1468), .A(n1463), .ZN(n122) );
  OAI21_X1 U520 ( .B1(N566), .B2(n1468), .A(n1463), .ZN(n367) );
  OAI21_X1 U521 ( .B1(N582), .B2(n1467), .A(n1464), .ZN(n205) );
  OAI21_X1 U522 ( .B1(N570), .B2(n1468), .A(n1463), .ZN(n325) );
  OAI21_X1 U523 ( .B1(N573), .B2(n1469), .A(n1464), .ZN(n296) );
  OAI21_X1 U524 ( .B1(N574), .B2(n1469), .A(n1464), .ZN(n288) );
  OAI21_X1 U525 ( .B1(DATA2[2]), .B2(n1467), .A(n453), .ZN(n467) );
  OAI21_X1 U526 ( .B1(DATA2[1]), .B2(n1467), .A(n453), .ZN(n474) );
  BUF_X1 U527 ( .A(n128), .Z(n1494) );
  OAI21_X1 U528 ( .B1(N555), .B2(n1467), .A(n1464), .ZN(n489) );
  INV_X1 U529 ( .A(n151), .ZN(n1610) );
  BUF_X1 U530 ( .A(N587), .Z(n1506) );
  BUF_X1 U531 ( .A(N587), .Z(n1507) );
  BUF_X1 U532 ( .A(N587), .Z(n1508) );
  INV_X1 U533 ( .A(DATA2[7]), .ZN(n1583) );
  INV_X1 U534 ( .A(DATA2[29]), .ZN(n1605) );
  INV_X1 U545 ( .A(DATA2[30]), .ZN(n1606) );
  INV_X1 U546 ( .A(DATA2[9]), .ZN(n1585) );
  INV_X1 U547 ( .A(DATA2[13]), .ZN(n1589) );
  INV_X1 U548 ( .A(DATA2[17]), .ZN(n1593) );
  INV_X1 U549 ( .A(DATA2[21]), .ZN(n1597) );
  INV_X1 U550 ( .A(DATA2[23]), .ZN(n1599) );
  INV_X1 U551 ( .A(DATA2[25]), .ZN(n1601) );
  INV_X1 U552 ( .A(DATA2[8]), .ZN(n1584) );
  INV_X1 U553 ( .A(DATA2[16]), .ZN(n1592) );
  INV_X1 U554 ( .A(DATA2[24]), .ZN(n1600) );
  INV_X1 U555 ( .A(DATA2[12]), .ZN(n1588) );
  INV_X1 U556 ( .A(DATA2[20]), .ZN(n1596) );
  INV_X1 U557 ( .A(DATA2[10]), .ZN(n1586) );
  INV_X1 U558 ( .A(DATA2[14]), .ZN(n1590) );
  INV_X1 U559 ( .A(DATA2[22]), .ZN(n1598) );
  INV_X1 U560 ( .A(DATA2[26]), .ZN(n1602) );
  NAND4_X1 U561 ( .A1(n485), .A2(n486), .A3(n487), .A4(n488), .ZN(N588) );
  AOI221_X1 U562 ( .B1(n380), .B2(n283), .C1(n332), .C2(n319), .A(n1529), .ZN(
        n486) );
  AOI221_X1 U563 ( .B1(DATA2[0]), .B2(n489), .C1(FUNC[3]), .C2(n490), .A(n491), 
        .ZN(n488) );
  AOI222_X1 U564 ( .A1(N389), .A2(n1482), .B1(n308), .B2(n361), .C1(N421), 
        .C2(n1485), .ZN(n485) );
  NAND2_X1 U565 ( .A1(N549), .A2(FUNC[0]), .ZN(n492) );
  NOR3_X1 U566 ( .A1(n493), .A2(FUNC[2]), .A3(n1609), .ZN(n138) );
  NOR3_X1 U567 ( .A1(FUNC[0]), .A2(FUNC[2]), .A3(n493), .ZN(n139) );
  AOI22_X1 U568 ( .A1(N550), .A2(n1609), .B1(N551), .B2(FUNC[0]), .ZN(n499) );
  AOI22_X1 U569 ( .A1(N552), .A2(n1609), .B1(N553), .B2(FUNC[0]), .ZN(n498) );
  NAND2_X1 U570 ( .A1(n504), .A2(FUNC[0]), .ZN(N587) );
  NAND2_X1 U571 ( .A1(n495), .A2(n496), .ZN(n490) );
  NAND2_X1 U572 ( .A1(n497), .A2(n1612), .ZN(n495) );
  NAND4_X1 U573 ( .A1(N554), .A2(FUNC[2]), .A3(n1609), .A4(n1611), .ZN(n496)
         );
  OAI22_X1 U574 ( .A1(n498), .A2(n1611), .B1(FUNC[1]), .B2(n499), .ZN(n497) );
  INV_X1 U575 ( .A(FUNC[0]), .ZN(n1609) );
  INV_X1 U576 ( .A(FUNC[2]), .ZN(n1612) );
  OR2_X1 U577 ( .A1(n1611), .A2(FUNC[3]), .ZN(n493) );
  INV_X1 U578 ( .A(FUNC[1]), .ZN(n1611) );
  OR3_X1 U579 ( .A1(FUNC[1]), .A2(FUNC[3]), .A3(n1612), .ZN(n128) );
  NOR3_X1 U580 ( .A1(FUNC[2]), .A2(FUNC[3]), .A3(FUNC[1]), .ZN(n317) );
  AND3_X1 U581 ( .A1(FUNC[2]), .A2(FUNC[1]), .A3(FUNC[3]), .ZN(n504) );
  INV_X1 U582 ( .A(n1454), .ZN(n1474) );
  INV_X1 U583 ( .A(n1454), .ZN(n1475) );
  INV_X1 U584 ( .A(n1454), .ZN(n1476) );
  INV_X1 U585 ( .A(n1453), .ZN(n1479) );
  INV_X1 U586 ( .A(n164), .ZN(n1481) );
  INV_X1 U587 ( .A(n129), .ZN(n1491) );
  INV_X1 U588 ( .A(n1502), .ZN(n1501) );
  INV_X1 U589 ( .A(n125), .ZN(n1502) );
endmodule


module FD_106 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_105 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_104 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_103 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_102 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_101 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_100 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_99 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_98 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_97 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_96 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_95 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_94 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_93 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_92 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_91 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_90 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_89 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_88 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_87 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_86 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_85 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_84 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_83 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_82 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_81 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_80 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_79 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_78 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_77 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_76 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_75 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_3 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_106 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_105 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_104 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_103 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_102 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_101 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_100 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_99 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_98 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_97 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_96 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_95 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_94 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_93 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_92 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_91 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_90 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_89 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_88 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_87 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_86 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_85 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_84 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_83 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_82 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_81 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_80 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_79 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_78 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_77 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_76 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_75 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FD_74 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_73 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_72 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_71 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_70 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_69 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_68 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_67 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_66 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_65 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_64 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_63 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_62 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_61 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_60 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_59 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_58 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_57 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_56 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_55 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_54 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_53 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_52 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_51 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_50 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_49 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_48 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_47 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_46 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_45 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_44 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_43 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_2 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_74 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_73 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_72 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_71 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_70 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_69 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_68 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_67 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_66 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_65 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_64 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_63 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_62 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_61 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_60 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_59 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_58 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_57 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_56 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_55 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_54 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_53 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_52 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_51 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_50 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_49 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_48 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_47 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_46 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_45 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_44 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_43 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module FD_42 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_41 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_40 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_39 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_38 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT5_2 ( D, CK, RESET, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  FD_42 UFD_0 ( .D(D[0]), .CK(CK), .RESET(RESET), .Q(Q[0]) );
  FD_41 UFD_1 ( .D(D[1]), .CK(CK), .RESET(RESET), .Q(Q[1]) );
  FD_40 UFD_2 ( .D(D[2]), .CK(CK), .RESET(RESET), .Q(Q[2]) );
  FD_39 UFD_3 ( .D(D[3]), .CK(CK), .RESET(RESET), .Q(Q[3]) );
  FD_38 UFD_4 ( .D(D[4]), .CK(CK), .RESET(RESET), .Q(Q[4]) );
endmodule


module EXECUTION_STAGE_numbit32 ( alu_forwarding_one, mem_forwarding_one, 
        alu_forwarding_two, mem_forwarding_two, alu_forwarding_value, 
        mem_forwarding_value, npc_in, a_reg_in, b_reg_in, imm_reg_in, 
        rd_reg_in, mux_one_control, mux_two_control, alu_control, clk, reset, 
        execution_stage_out, b_reg_out, rd_reg_out );
  input [31:0] alu_forwarding_value;
  input [31:0] mem_forwarding_value;
  input [31:0] npc_in;
  input [31:0] a_reg_in;
  input [31:0] b_reg_in;
  input [31:0] imm_reg_in;
  input [4:0] rd_reg_in;
  input [3:0] alu_control;
  output [31:0] execution_stage_out;
  output [31:0] b_reg_out;
  output [4:0] rd_reg_out;
  input alu_forwarding_one, mem_forwarding_one, alu_forwarding_two,
         mem_forwarding_two, mux_one_control, mux_two_control, clk, reset;

  wire   [31:0] mux_one_out_rf;
  wire   [31:0] mux_one_out_mem_forwarding;
  wire   [31:0] mux_one_out_alu_forwarding;
  wire   [31:0] mux_two_out_rf;
  wire   [31:0] mux_two_out_mem_forwarding;
  wire   [31:0] mux_two_out_alu_forwarding;
  wire   [31:0] alu_out;

  MUX21_GENERIC_NBIT32_0 MUX_ONE_RF ( .A(npc_in), .B(a_reg_in), .SEL(
        mux_one_control), .Y(mux_one_out_rf) );
  MUX21_GENERIC_NBIT32_6 MUX_ONE_MEM ( .A(mux_one_out_rf), .B(
        mem_forwarding_value), .SEL(mem_forwarding_one), .Y(
        mux_one_out_mem_forwarding) );
  MUX21_GENERIC_NBIT32_5 MUX_ONE_ALU ( .A(mux_one_out_mem_forwarding), .B(
        alu_forwarding_value), .SEL(alu_forwarding_one), .Y(
        mux_one_out_alu_forwarding) );
  MUX21_GENERIC_NBIT32_4 MUX_TWO_RF ( .A(b_reg_in), .B(imm_reg_in), .SEL(
        mux_two_control), .Y(mux_two_out_rf) );
  MUX21_GENERIC_NBIT32_3 MUX_TWO_MEM ( .A(mux_two_out_rf), .B(
        mem_forwarding_value), .SEL(mem_forwarding_two), .Y(
        mux_two_out_mem_forwarding) );
  MUX21_GENERIC_NBIT32_2 MUX_TWO_ALU ( .A(mux_two_out_mem_forwarding), .B(
        alu_forwarding_value), .SEL(alu_forwarding_two), .Y(
        mux_two_out_alu_forwarding) );
  ALU_BEHAVIORAL_NBIT32 ALU ( .FUNC(alu_control), .DATA1(
        mux_one_out_alu_forwarding), .DATA2(mux_two_out_alu_forwarding), 
        .OUTALU(alu_out) );
  REGISTER_GENERIC_NBIT32_3 REG1 ( .D(alu_out), .CK(clk), .RESET(reset), .Q(
        execution_stage_out) );
  REGISTER_GENERIC_NBIT32_2 REG3 ( .D(b_reg_in), .CK(clk), .RESET(reset), .Q(
        b_reg_out) );
  REGISTER_GENERIC_NBIT5_2 REG4 ( .D(rd_reg_in), .CK(clk), .RESET(reset), .Q(
        rd_reg_out) );
endmodule


module FD_37 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_36 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_35 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_34 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_33 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT5_1 ( D, CK, RESET, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET;


  FD_37 UFD_0 ( .D(D[0]), .CK(CK), .RESET(RESET), .Q(Q[0]) );
  FD_36 UFD_1 ( .D(D[1]), .CK(CK), .RESET(RESET), .Q(Q[1]) );
  FD_35 UFD_2 ( .D(D[2]), .CK(CK), .RESET(RESET), .Q(Q[2]) );
  FD_34 UFD_3 ( .D(D[3]), .CK(CK), .RESET(RESET), .Q(Q[3]) );
  FD_33 UFD_4 ( .D(D[4]), .CK(CK), .RESET(RESET), .Q(Q[4]) );
endmodule


module FD_32 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_31 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_30 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_29 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_28 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_27 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_26 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_25 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_24 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_23 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_22 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_21 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_20 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_19 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_18 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_17 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_16 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_15 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_14 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_13 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_12 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_11 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_10 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_9 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_8 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_7 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_6 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_5 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_4 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_3 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_2 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module FD_1 ( D, CK, RESET, Q );
  input D, CK, RESET;
  output Q;
  wire   N3, n7;

  DFF_X1 Q_reg ( .D(N3), .CK(CK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n7), .ZN(N3) );
  INV_X1 U4 ( .A(D), .ZN(n7) );
endmodule


module REGISTER_GENERIC_NBIT32_1 ( D, CK, RESET, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET;
  wire   n19, n20, n21;

  FD_32 UFD_0 ( .D(D[0]), .CK(CK), .RESET(n19), .Q(Q[0]) );
  FD_31 UFD_1 ( .D(D[1]), .CK(CK), .RESET(n19), .Q(Q[1]) );
  FD_30 UFD_2 ( .D(D[2]), .CK(CK), .RESET(n19), .Q(Q[2]) );
  FD_29 UFD_3 ( .D(D[3]), .CK(CK), .RESET(n19), .Q(Q[3]) );
  FD_28 UFD_4 ( .D(D[4]), .CK(CK), .RESET(n19), .Q(Q[4]) );
  FD_27 UFD_5 ( .D(D[5]), .CK(CK), .RESET(n19), .Q(Q[5]) );
  FD_26 UFD_6 ( .D(D[6]), .CK(CK), .RESET(n19), .Q(Q[6]) );
  FD_25 UFD_7 ( .D(D[7]), .CK(CK), .RESET(n19), .Q(Q[7]) );
  FD_24 UFD_8 ( .D(D[8]), .CK(CK), .RESET(n19), .Q(Q[8]) );
  FD_23 UFD_9 ( .D(D[9]), .CK(CK), .RESET(n19), .Q(Q[9]) );
  FD_22 UFD_10 ( .D(D[10]), .CK(CK), .RESET(n19), .Q(Q[10]) );
  FD_21 UFD_11 ( .D(D[11]), .CK(CK), .RESET(n19), .Q(Q[11]) );
  FD_20 UFD_12 ( .D(D[12]), .CK(CK), .RESET(n20), .Q(Q[12]) );
  FD_19 UFD_13 ( .D(D[13]), .CK(CK), .RESET(n20), .Q(Q[13]) );
  FD_18 UFD_14 ( .D(D[14]), .CK(CK), .RESET(n20), .Q(Q[14]) );
  FD_17 UFD_15 ( .D(D[15]), .CK(CK), .RESET(n20), .Q(Q[15]) );
  FD_16 UFD_16 ( .D(D[16]), .CK(CK), .RESET(n20), .Q(Q[16]) );
  FD_15 UFD_17 ( .D(D[17]), .CK(CK), .RESET(n20), .Q(Q[17]) );
  FD_14 UFD_18 ( .D(D[18]), .CK(CK), .RESET(n20), .Q(Q[18]) );
  FD_13 UFD_19 ( .D(D[19]), .CK(CK), .RESET(n20), .Q(Q[19]) );
  FD_12 UFD_20 ( .D(D[20]), .CK(CK), .RESET(n20), .Q(Q[20]) );
  FD_11 UFD_21 ( .D(D[21]), .CK(CK), .RESET(n20), .Q(Q[21]) );
  FD_10 UFD_22 ( .D(D[22]), .CK(CK), .RESET(n20), .Q(Q[22]) );
  FD_9 UFD_23 ( .D(D[23]), .CK(CK), .RESET(n20), .Q(Q[23]) );
  FD_8 UFD_24 ( .D(D[24]), .CK(CK), .RESET(n21), .Q(Q[24]) );
  FD_7 UFD_25 ( .D(D[25]), .CK(CK), .RESET(n21), .Q(Q[25]) );
  FD_6 UFD_26 ( .D(D[26]), .CK(CK), .RESET(n21), .Q(Q[26]) );
  FD_5 UFD_27 ( .D(D[27]), .CK(CK), .RESET(n21), .Q(Q[27]) );
  FD_4 UFD_28 ( .D(D[28]), .CK(CK), .RESET(n21), .Q(Q[28]) );
  FD_3 UFD_29 ( .D(D[29]), .CK(CK), .RESET(n21), .Q(Q[29]) );
  FD_2 UFD_30 ( .D(D[30]), .CK(CK), .RESET(n21), .Q(Q[30]) );
  FD_1 UFD_31 ( .D(D[31]), .CK(CK), .RESET(n21), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RESET), .Z(n19) );
  BUF_X1 U2 ( .A(RESET), .Z(n20) );
  BUF_X1 U3 ( .A(RESET), .Z(n21) );
endmodule


module MEMORY_STAGE_numbit32 ( alu_in, rd_reg_in, reset, clk, to_mem_stage_reg, 
        rd_reg_out, memory_stage_out, alu_out );
  input [31:0] alu_in;
  input [4:0] rd_reg_in;
  input [31:0] to_mem_stage_reg;
  output [4:0] rd_reg_out;
  output [31:0] memory_stage_out;
  output [31:0] alu_out;
  input reset, clk;

  assign memory_stage_out[31] = to_mem_stage_reg[31];
  assign memory_stage_out[30] = to_mem_stage_reg[30];
  assign memory_stage_out[29] = to_mem_stage_reg[29];
  assign memory_stage_out[28] = to_mem_stage_reg[28];
  assign memory_stage_out[27] = to_mem_stage_reg[27];
  assign memory_stage_out[26] = to_mem_stage_reg[26];
  assign memory_stage_out[25] = to_mem_stage_reg[25];
  assign memory_stage_out[24] = to_mem_stage_reg[24];
  assign memory_stage_out[23] = to_mem_stage_reg[23];
  assign memory_stage_out[22] = to_mem_stage_reg[22];
  assign memory_stage_out[21] = to_mem_stage_reg[21];
  assign memory_stage_out[20] = to_mem_stage_reg[20];
  assign memory_stage_out[19] = to_mem_stage_reg[19];
  assign memory_stage_out[18] = to_mem_stage_reg[18];
  assign memory_stage_out[17] = to_mem_stage_reg[17];
  assign memory_stage_out[16] = to_mem_stage_reg[16];
  assign memory_stage_out[15] = to_mem_stage_reg[15];
  assign memory_stage_out[14] = to_mem_stage_reg[14];
  assign memory_stage_out[13] = to_mem_stage_reg[13];
  assign memory_stage_out[12] = to_mem_stage_reg[12];
  assign memory_stage_out[11] = to_mem_stage_reg[11];
  assign memory_stage_out[10] = to_mem_stage_reg[10];
  assign memory_stage_out[9] = to_mem_stage_reg[9];
  assign memory_stage_out[8] = to_mem_stage_reg[8];
  assign memory_stage_out[7] = to_mem_stage_reg[7];
  assign memory_stage_out[6] = to_mem_stage_reg[6];
  assign memory_stage_out[5] = to_mem_stage_reg[5];
  assign memory_stage_out[4] = to_mem_stage_reg[4];
  assign memory_stage_out[3] = to_mem_stage_reg[3];
  assign memory_stage_out[2] = to_mem_stage_reg[2];
  assign memory_stage_out[1] = to_mem_stage_reg[1];
  assign memory_stage_out[0] = to_mem_stage_reg[0];

  REGISTER_GENERIC_NBIT5_1 RDREG ( .D(rd_reg_in), .CK(clk), .RESET(reset), .Q(
        rd_reg_out) );
  REGISTER_GENERIC_NBIT32_1 REGALU ( .D(alu_in), .CK(clk), .RESET(reset), .Q(
        alu_out) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;

  wire   [31:0] SEL_INV;
  wire   [31:0] NAND_ONE_OUT;
  wire   [31:0] NAND_TWO_OUT;

  IV_37 UIV_0 ( .A(SEL), .Y(SEL_INV[0]) );
  ND2_111 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_110 UND2_0 ( .A(B[0]), .B(SEL), .Y(NAND_TWO_OUT[0]) );
  ND2_109 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_36 UIV_1 ( .A(SEL), .Y(SEL_INV[1]) );
  ND2_108 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_107 UND2_1 ( .A(B[1]), .B(SEL), .Y(NAND_TWO_OUT[1]) );
  ND2_106 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_35 UIV_2 ( .A(SEL), .Y(SEL_INV[2]) );
  ND2_105 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_104 UND2_2 ( .A(B[2]), .B(SEL), .Y(NAND_TWO_OUT[2]) );
  ND2_103 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_34 UIV_3 ( .A(SEL), .Y(SEL_INV[3]) );
  ND2_102 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_101 UND2_3 ( .A(B[3]), .B(SEL), .Y(NAND_TWO_OUT[3]) );
  ND2_100 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_33 UIV_4 ( .A(SEL), .Y(SEL_INV[4]) );
  ND2_99 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_98 UND2_4 ( .A(B[4]), .B(SEL), .Y(NAND_TWO_OUT[4]) );
  ND2_97 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
  IV_32 UIV_5 ( .A(SEL), .Y(SEL_INV[5]) );
  ND2_96 UND1_5 ( .A(A[5]), .B(SEL_INV[5]), .Y(NAND_ONE_OUT[5]) );
  ND2_95 UND2_5 ( .A(B[5]), .B(SEL), .Y(NAND_TWO_OUT[5]) );
  ND2_94 UND3_5 ( .A(NAND_ONE_OUT[5]), .B(NAND_TWO_OUT[5]), .Y(Y[5]) );
  IV_31 UIV_6 ( .A(SEL), .Y(SEL_INV[6]) );
  ND2_93 UND1_6 ( .A(A[6]), .B(SEL_INV[6]), .Y(NAND_ONE_OUT[6]) );
  ND2_92 UND2_6 ( .A(B[6]), .B(SEL), .Y(NAND_TWO_OUT[6]) );
  ND2_91 UND3_6 ( .A(NAND_ONE_OUT[6]), .B(NAND_TWO_OUT[6]), .Y(Y[6]) );
  IV_30 UIV_7 ( .A(SEL), .Y(SEL_INV[7]) );
  ND2_90 UND1_7 ( .A(A[7]), .B(SEL_INV[7]), .Y(NAND_ONE_OUT[7]) );
  ND2_89 UND2_7 ( .A(B[7]), .B(SEL), .Y(NAND_TWO_OUT[7]) );
  ND2_88 UND3_7 ( .A(NAND_ONE_OUT[7]), .B(NAND_TWO_OUT[7]), .Y(Y[7]) );
  IV_29 UIV_8 ( .A(SEL), .Y(SEL_INV[8]) );
  ND2_87 UND1_8 ( .A(A[8]), .B(SEL_INV[8]), .Y(NAND_ONE_OUT[8]) );
  ND2_86 UND2_8 ( .A(B[8]), .B(SEL), .Y(NAND_TWO_OUT[8]) );
  ND2_85 UND3_8 ( .A(NAND_ONE_OUT[8]), .B(NAND_TWO_OUT[8]), .Y(Y[8]) );
  IV_28 UIV_9 ( .A(SEL), .Y(SEL_INV[9]) );
  ND2_84 UND1_9 ( .A(A[9]), .B(SEL_INV[9]), .Y(NAND_ONE_OUT[9]) );
  ND2_83 UND2_9 ( .A(B[9]), .B(SEL), .Y(NAND_TWO_OUT[9]) );
  ND2_82 UND3_9 ( .A(NAND_ONE_OUT[9]), .B(NAND_TWO_OUT[9]), .Y(Y[9]) );
  IV_27 UIV_10 ( .A(SEL), .Y(SEL_INV[10]) );
  ND2_81 UND1_10 ( .A(A[10]), .B(SEL_INV[10]), .Y(NAND_ONE_OUT[10]) );
  ND2_80 UND2_10 ( .A(B[10]), .B(SEL), .Y(NAND_TWO_OUT[10]) );
  ND2_79 UND3_10 ( .A(NAND_ONE_OUT[10]), .B(NAND_TWO_OUT[10]), .Y(Y[10]) );
  IV_26 UIV_11 ( .A(SEL), .Y(SEL_INV[11]) );
  ND2_78 UND1_11 ( .A(A[11]), .B(SEL_INV[11]), .Y(NAND_ONE_OUT[11]) );
  ND2_77 UND2_11 ( .A(B[11]), .B(SEL), .Y(NAND_TWO_OUT[11]) );
  ND2_76 UND3_11 ( .A(NAND_ONE_OUT[11]), .B(NAND_TWO_OUT[11]), .Y(Y[11]) );
  IV_25 UIV_12 ( .A(SEL), .Y(SEL_INV[12]) );
  ND2_75 UND1_12 ( .A(A[12]), .B(SEL_INV[12]), .Y(NAND_ONE_OUT[12]) );
  ND2_74 UND2_12 ( .A(B[12]), .B(SEL), .Y(NAND_TWO_OUT[12]) );
  ND2_73 UND3_12 ( .A(NAND_ONE_OUT[12]), .B(NAND_TWO_OUT[12]), .Y(Y[12]) );
  IV_24 UIV_13 ( .A(SEL), .Y(SEL_INV[13]) );
  ND2_72 UND1_13 ( .A(A[13]), .B(SEL_INV[13]), .Y(NAND_ONE_OUT[13]) );
  ND2_71 UND2_13 ( .A(B[13]), .B(SEL), .Y(NAND_TWO_OUT[13]) );
  ND2_70 UND3_13 ( .A(NAND_ONE_OUT[13]), .B(NAND_TWO_OUT[13]), .Y(Y[13]) );
  IV_23 UIV_14 ( .A(SEL), .Y(SEL_INV[14]) );
  ND2_69 UND1_14 ( .A(A[14]), .B(SEL_INV[14]), .Y(NAND_ONE_OUT[14]) );
  ND2_68 UND2_14 ( .A(B[14]), .B(SEL), .Y(NAND_TWO_OUT[14]) );
  ND2_67 UND3_14 ( .A(NAND_ONE_OUT[14]), .B(NAND_TWO_OUT[14]), .Y(Y[14]) );
  IV_22 UIV_15 ( .A(SEL), .Y(SEL_INV[15]) );
  ND2_66 UND1_15 ( .A(A[15]), .B(SEL_INV[15]), .Y(NAND_ONE_OUT[15]) );
  ND2_65 UND2_15 ( .A(B[15]), .B(SEL), .Y(NAND_TWO_OUT[15]) );
  ND2_64 UND3_15 ( .A(NAND_ONE_OUT[15]), .B(NAND_TWO_OUT[15]), .Y(Y[15]) );
  IV_21 UIV_16 ( .A(SEL), .Y(SEL_INV[16]) );
  ND2_63 UND1_16 ( .A(A[16]), .B(SEL_INV[16]), .Y(NAND_ONE_OUT[16]) );
  ND2_62 UND2_16 ( .A(B[16]), .B(SEL), .Y(NAND_TWO_OUT[16]) );
  ND2_61 UND3_16 ( .A(NAND_ONE_OUT[16]), .B(NAND_TWO_OUT[16]), .Y(Y[16]) );
  IV_20 UIV_17 ( .A(SEL), .Y(SEL_INV[17]) );
  ND2_60 UND1_17 ( .A(A[17]), .B(SEL_INV[17]), .Y(NAND_ONE_OUT[17]) );
  ND2_59 UND2_17 ( .A(B[17]), .B(SEL), .Y(NAND_TWO_OUT[17]) );
  ND2_58 UND3_17 ( .A(NAND_ONE_OUT[17]), .B(NAND_TWO_OUT[17]), .Y(Y[17]) );
  IV_19 UIV_18 ( .A(SEL), .Y(SEL_INV[18]) );
  ND2_57 UND1_18 ( .A(A[18]), .B(SEL_INV[18]), .Y(NAND_ONE_OUT[18]) );
  ND2_56 UND2_18 ( .A(B[18]), .B(SEL), .Y(NAND_TWO_OUT[18]) );
  ND2_55 UND3_18 ( .A(NAND_ONE_OUT[18]), .B(NAND_TWO_OUT[18]), .Y(Y[18]) );
  IV_18 UIV_19 ( .A(SEL), .Y(SEL_INV[19]) );
  ND2_54 UND1_19 ( .A(A[19]), .B(SEL_INV[19]), .Y(NAND_ONE_OUT[19]) );
  ND2_53 UND2_19 ( .A(B[19]), .B(SEL), .Y(NAND_TWO_OUT[19]) );
  ND2_52 UND3_19 ( .A(NAND_ONE_OUT[19]), .B(NAND_TWO_OUT[19]), .Y(Y[19]) );
  IV_17 UIV_20 ( .A(SEL), .Y(SEL_INV[20]) );
  ND2_51 UND1_20 ( .A(A[20]), .B(SEL_INV[20]), .Y(NAND_ONE_OUT[20]) );
  ND2_50 UND2_20 ( .A(B[20]), .B(SEL), .Y(NAND_TWO_OUT[20]) );
  ND2_49 UND3_20 ( .A(NAND_ONE_OUT[20]), .B(NAND_TWO_OUT[20]), .Y(Y[20]) );
  IV_16 UIV_21 ( .A(SEL), .Y(SEL_INV[21]) );
  ND2_48 UND1_21 ( .A(A[21]), .B(SEL_INV[21]), .Y(NAND_ONE_OUT[21]) );
  ND2_47 UND2_21 ( .A(B[21]), .B(SEL), .Y(NAND_TWO_OUT[21]) );
  ND2_46 UND3_21 ( .A(NAND_ONE_OUT[21]), .B(NAND_TWO_OUT[21]), .Y(Y[21]) );
  IV_15 UIV_22 ( .A(SEL), .Y(SEL_INV[22]) );
  ND2_45 UND1_22 ( .A(A[22]), .B(SEL_INV[22]), .Y(NAND_ONE_OUT[22]) );
  ND2_44 UND2_22 ( .A(B[22]), .B(SEL), .Y(NAND_TWO_OUT[22]) );
  ND2_43 UND3_22 ( .A(NAND_ONE_OUT[22]), .B(NAND_TWO_OUT[22]), .Y(Y[22]) );
  IV_14 UIV_23 ( .A(SEL), .Y(SEL_INV[23]) );
  ND2_42 UND1_23 ( .A(A[23]), .B(SEL_INV[23]), .Y(NAND_ONE_OUT[23]) );
  ND2_41 UND2_23 ( .A(B[23]), .B(SEL), .Y(NAND_TWO_OUT[23]) );
  ND2_40 UND3_23 ( .A(NAND_ONE_OUT[23]), .B(NAND_TWO_OUT[23]), .Y(Y[23]) );
  IV_13 UIV_24 ( .A(SEL), .Y(SEL_INV[24]) );
  ND2_39 UND1_24 ( .A(A[24]), .B(SEL_INV[24]), .Y(NAND_ONE_OUT[24]) );
  ND2_38 UND2_24 ( .A(B[24]), .B(SEL), .Y(NAND_TWO_OUT[24]) );
  ND2_37 UND3_24 ( .A(NAND_ONE_OUT[24]), .B(NAND_TWO_OUT[24]), .Y(Y[24]) );
  IV_12 UIV_25 ( .A(SEL), .Y(SEL_INV[25]) );
  ND2_36 UND1_25 ( .A(A[25]), .B(SEL_INV[25]), .Y(NAND_ONE_OUT[25]) );
  ND2_35 UND2_25 ( .A(B[25]), .B(SEL), .Y(NAND_TWO_OUT[25]) );
  ND2_34 UND3_25 ( .A(NAND_ONE_OUT[25]), .B(NAND_TWO_OUT[25]), .Y(Y[25]) );
  IV_11 UIV_26 ( .A(SEL), .Y(SEL_INV[26]) );
  ND2_33 UND1_26 ( .A(A[26]), .B(SEL_INV[26]), .Y(NAND_ONE_OUT[26]) );
  ND2_32 UND2_26 ( .A(B[26]), .B(SEL), .Y(NAND_TWO_OUT[26]) );
  ND2_31 UND3_26 ( .A(NAND_ONE_OUT[26]), .B(NAND_TWO_OUT[26]), .Y(Y[26]) );
  IV_10 UIV_27 ( .A(SEL), .Y(SEL_INV[27]) );
  ND2_30 UND1_27 ( .A(A[27]), .B(SEL_INV[27]), .Y(NAND_ONE_OUT[27]) );
  ND2_29 UND2_27 ( .A(B[27]), .B(SEL), .Y(NAND_TWO_OUT[27]) );
  ND2_28 UND3_27 ( .A(NAND_ONE_OUT[27]), .B(NAND_TWO_OUT[27]), .Y(Y[27]) );
  IV_9 UIV_28 ( .A(SEL), .Y(SEL_INV[28]) );
  ND2_27 UND1_28 ( .A(A[28]), .B(SEL_INV[28]), .Y(NAND_ONE_OUT[28]) );
  ND2_26 UND2_28 ( .A(B[28]), .B(SEL), .Y(NAND_TWO_OUT[28]) );
  ND2_25 UND3_28 ( .A(NAND_ONE_OUT[28]), .B(NAND_TWO_OUT[28]), .Y(Y[28]) );
  IV_8 UIV_29 ( .A(SEL), .Y(SEL_INV[29]) );
  ND2_24 UND1_29 ( .A(A[29]), .B(SEL_INV[29]), .Y(NAND_ONE_OUT[29]) );
  ND2_23 UND2_29 ( .A(B[29]), .B(SEL), .Y(NAND_TWO_OUT[29]) );
  ND2_22 UND3_29 ( .A(NAND_ONE_OUT[29]), .B(NAND_TWO_OUT[29]), .Y(Y[29]) );
  IV_7 UIV_30 ( .A(SEL), .Y(SEL_INV[30]) );
  ND2_21 UND1_30 ( .A(A[30]), .B(SEL_INV[30]), .Y(NAND_ONE_OUT[30]) );
  ND2_20 UND2_30 ( .A(B[30]), .B(SEL), .Y(NAND_TWO_OUT[30]) );
  ND2_19 UND3_30 ( .A(NAND_ONE_OUT[30]), .B(NAND_TWO_OUT[30]), .Y(Y[30]) );
  IV_6 UIV_31 ( .A(SEL), .Y(SEL_INV[31]) );
  ND2_18 UND1_31 ( .A(A[31]), .B(SEL_INV[31]), .Y(NAND_ONE_OUT[31]) );
  ND2_17 UND2_31 ( .A(B[31]), .B(SEL), .Y(NAND_TWO_OUT[31]) );
  ND2_16 UND3_31 ( .A(NAND_ONE_OUT[31]), .B(NAND_TWO_OUT[31]), .Y(Y[31]) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT5 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;

  wire   [4:0] SEL_INV;
  wire   [4:0] NAND_ONE_OUT;
  wire   [4:0] NAND_TWO_OUT;

  IV_5 UIV_0 ( .A(SEL), .Y(SEL_INV[0]) );
  ND2_15 UND1_0 ( .A(A[0]), .B(SEL_INV[0]), .Y(NAND_ONE_OUT[0]) );
  ND2_14 UND2_0 ( .A(B[0]), .B(SEL), .Y(NAND_TWO_OUT[0]) );
  ND2_13 UND3_0 ( .A(NAND_ONE_OUT[0]), .B(NAND_TWO_OUT[0]), .Y(Y[0]) );
  IV_4 UIV_1 ( .A(SEL), .Y(SEL_INV[1]) );
  ND2_12 UND1_1 ( .A(A[1]), .B(SEL_INV[1]), .Y(NAND_ONE_OUT[1]) );
  ND2_11 UND2_1 ( .A(B[1]), .B(SEL), .Y(NAND_TWO_OUT[1]) );
  ND2_10 UND3_1 ( .A(NAND_ONE_OUT[1]), .B(NAND_TWO_OUT[1]), .Y(Y[1]) );
  IV_3 UIV_2 ( .A(SEL), .Y(SEL_INV[2]) );
  ND2_9 UND1_2 ( .A(A[2]), .B(SEL_INV[2]), .Y(NAND_ONE_OUT[2]) );
  ND2_8 UND2_2 ( .A(B[2]), .B(SEL), .Y(NAND_TWO_OUT[2]) );
  ND2_7 UND3_2 ( .A(NAND_ONE_OUT[2]), .B(NAND_TWO_OUT[2]), .Y(Y[2]) );
  IV_2 UIV_3 ( .A(SEL), .Y(SEL_INV[3]) );
  ND2_6 UND1_3 ( .A(A[3]), .B(SEL_INV[3]), .Y(NAND_ONE_OUT[3]) );
  ND2_5 UND2_3 ( .A(B[3]), .B(SEL), .Y(NAND_TWO_OUT[3]) );
  ND2_4 UND3_3 ( .A(NAND_ONE_OUT[3]), .B(NAND_TWO_OUT[3]), .Y(Y[3]) );
  IV_1 UIV_4 ( .A(SEL), .Y(SEL_INV[4]) );
  ND2_3 UND1_4 ( .A(A[4]), .B(SEL_INV[4]), .Y(NAND_ONE_OUT[4]) );
  ND2_2 UND2_4 ( .A(B[4]), .B(SEL), .Y(NAND_TWO_OUT[4]) );
  ND2_1 UND3_4 ( .A(NAND_ONE_OUT[4]), .B(NAND_TWO_OUT[4]), .Y(Y[4]) );
endmodule


module WRITE_BACK_STAGE_N32 ( LMD, ALUOUT, RD_IN, CONTROL, JAL_SEL, RD_OUT, 
        WB_OUT );
  input [31:0] LMD;
  input [31:0] ALUOUT;
  input [4:0] RD_IN;
  output [4:0] RD_OUT;
  output [31:0] WB_OUT;
  input CONTROL, JAL_SEL;


  MUX21_GENERIC_NBIT32_1 UMUX ( .A(LMD), .B(ALUOUT), .SEL(CONTROL), .Y(WB_OUT)
         );
  MUX21_GENERIC_NBIT5 JALMUX ( .A(RD_IN), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .SEL(JAL_SEL), .Y(RD_OUT) );
endmodule


module DATAPATH_numbit32 ( clk, reset, write_enable, mux_one_control, 
        mux_two_control, alu_control, to_ir, to_mem_stage_reg, wb_control, 
        jal_sel, to_iram, npc_out_if, npc_out_bpu, instruction_fetched, ir_out, 
        rd_out_id, npc_out_id, a_reg_out, b_reg_out, imm_reg_out, alu_out, 
        rd_out_ex, b_reg_out_ex, rd_out_mem, memory_stage_out, alu_out_mem, 
        wb_stage_out, rd_out_wb, alu_forwarding_one, mem_forwarding_one, 
        alu_forwarding_two, mem_forwarding_two, alu_forwarding_value, 
        mem_forwarding_value );
  input [3:0] alu_control;
  input [31:0] to_ir;
  input [31:0] to_mem_stage_reg;
  output [31:0] to_iram;
  output [31:0] npc_out_if;
  output [31:0] npc_out_bpu;
  output [31:0] instruction_fetched;
  output [31:0] ir_out;
  output [4:0] rd_out_id;
  output [31:0] npc_out_id;
  output [31:0] a_reg_out;
  output [31:0] b_reg_out;
  output [31:0] imm_reg_out;
  output [31:0] alu_out;
  output [4:0] rd_out_ex;
  output [31:0] b_reg_out_ex;
  output [4:0] rd_out_mem;
  output [31:0] memory_stage_out;
  output [31:0] alu_out_mem;
  output [31:0] wb_stage_out;
  output [4:0] rd_out_wb;
  output [31:0] alu_forwarding_value;
  output [31:0] mem_forwarding_value;
  input clk, reset, write_enable, mux_one_control, mux_two_control, wb_control,
         jal_sel;
  output alu_forwarding_one, mem_forwarding_one, alu_forwarding_two,
         mem_forwarding_two;
  wire   n4, n9;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign to_iram[31] = 1'b0;
  assign to_iram[30] = 1'b0;
  assign ir_out[22] = n4;
  assign alu_forwarding_value[31] = alu_out[31];
  assign alu_forwarding_value[30] = alu_out[30];
  assign alu_forwarding_value[29] = alu_out[29];
  assign alu_forwarding_value[28] = alu_out[28];
  assign alu_forwarding_value[27] = alu_out[27];
  assign alu_forwarding_value[26] = alu_out[26];
  assign alu_forwarding_value[25] = alu_out[25];
  assign alu_forwarding_value[24] = alu_out[24];
  assign alu_forwarding_value[23] = alu_out[23];
  assign alu_forwarding_value[22] = alu_out[22];
  assign alu_forwarding_value[21] = alu_out[21];
  assign alu_forwarding_value[20] = alu_out[20];
  assign alu_forwarding_value[19] = alu_out[19];
  assign alu_forwarding_value[18] = alu_out[18];
  assign alu_forwarding_value[17] = alu_out[17];
  assign alu_forwarding_value[16] = alu_out[16];
  assign alu_forwarding_value[15] = alu_out[15];
  assign alu_forwarding_value[14] = alu_out[14];
  assign alu_forwarding_value[13] = alu_out[13];
  assign alu_forwarding_value[12] = alu_out[12];
  assign alu_forwarding_value[11] = alu_out[11];
  assign alu_forwarding_value[10] = alu_out[10];
  assign alu_forwarding_value[9] = alu_out[9];
  assign alu_forwarding_value[8] = alu_out[8];
  assign alu_forwarding_value[7] = alu_out[7];
  assign alu_forwarding_value[6] = alu_out[6];
  assign alu_forwarding_value[5] = alu_out[5];
  assign alu_forwarding_value[4] = alu_out[4];
  assign alu_forwarding_value[3] = alu_out[3];
  assign alu_forwarding_value[2] = alu_out[2];
  assign alu_forwarding_value[1] = alu_out[1];
  assign alu_forwarding_value[0] = alu_out[0];
  assign mem_forwarding_value[31] = alu_out_mem[31];
  assign mem_forwarding_value[30] = alu_out_mem[30];
  assign mem_forwarding_value[29] = alu_out_mem[29];
  assign mem_forwarding_value[28] = alu_out_mem[28];
  assign mem_forwarding_value[27] = alu_out_mem[27];
  assign mem_forwarding_value[26] = alu_out_mem[26];
  assign mem_forwarding_value[25] = alu_out_mem[25];
  assign mem_forwarding_value[24] = alu_out_mem[24];
  assign mem_forwarding_value[23] = alu_out_mem[23];
  assign mem_forwarding_value[22] = alu_out_mem[22];
  assign mem_forwarding_value[21] = alu_out_mem[21];
  assign mem_forwarding_value[20] = alu_out_mem[20];
  assign mem_forwarding_value[19] = alu_out_mem[19];
  assign mem_forwarding_value[18] = alu_out_mem[18];
  assign mem_forwarding_value[17] = alu_out_mem[17];
  assign mem_forwarding_value[16] = alu_out_mem[16];
  assign mem_forwarding_value[15] = alu_out_mem[15];
  assign mem_forwarding_value[14] = alu_out_mem[14];
  assign mem_forwarding_value[13] = alu_out_mem[13];
  assign mem_forwarding_value[12] = alu_out_mem[12];
  assign mem_forwarding_value[11] = alu_out_mem[11];
  assign mem_forwarding_value[10] = alu_out_mem[10];
  assign mem_forwarding_value[9] = alu_out_mem[9];
  assign mem_forwarding_value[8] = alu_out_mem[8];
  assign mem_forwarding_value[7] = alu_out_mem[7];
  assign mem_forwarding_value[6] = alu_out_mem[6];
  assign mem_forwarding_value[5] = alu_out_mem[5];
  assign mem_forwarding_value[4] = alu_out_mem[4];
  assign mem_forwarding_value[3] = alu_out_mem[3];
  assign mem_forwarding_value[2] = alu_out_mem[2];
  assign mem_forwarding_value[1] = alu_out_mem[1];
  assign mem_forwarding_value[0] = alu_out_mem[0];

  FETCH_STAGE_numbit32 FETCH ( .program_counter(npc_out_bpu), .to_IR(to_ir), 
        .clk(clk), .reset(n9), .to_IRAM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, to_iram[29:0]}), .npc_out(npc_out_if), 
        .instruction_reg_out({ir_out[31:23], n4, ir_out[21:0]}), 
        .instruction_fetched(instruction_fetched) );
  DECODE_STAGE_numbit32 DECODE ( .IR_IN({ir_out[31:23], n4, ir_out[21:0]}), 
        .WB_STAGE_IN(wb_stage_out), .NPC_IN(npc_out_if), .RD_IN(rd_out_wb), 
        .CLK(clk), .RESET(n9), .WRITE_ENABLE(write_enable), 
        .INSTRUCTION_FETCHED(instruction_fetched), .NPC_OUT_BPU(npc_out_bpu), 
        .RD_OUT(rd_out_id), .NPC_OUT(npc_out_id), .A_REG_OUT(a_reg_out), 
        .B_REG_OUT(b_reg_out), .IMM_REG_OUT(imm_reg_out), .alu_forwarding_one(
        alu_forwarding_one), .mem_forwarding_one(mem_forwarding_one), 
        .alu_forwarding_two(alu_forwarding_two), .mem_forwarding_two(
        mem_forwarding_two) );
  EXECUTION_STAGE_numbit32 EXECUTE ( .alu_forwarding_one(alu_forwarding_one), 
        .mem_forwarding_one(mem_forwarding_one), .alu_forwarding_two(
        alu_forwarding_two), .mem_forwarding_two(mem_forwarding_two), 
        .alu_forwarding_value(alu_out), .mem_forwarding_value(alu_out_mem), 
        .npc_in(npc_out_id), .a_reg_in(a_reg_out), .b_reg_in(b_reg_out), 
        .imm_reg_in(imm_reg_out), .rd_reg_in(rd_out_id), .mux_one_control(
        mux_one_control), .mux_two_control(mux_two_control), .alu_control(
        alu_control), .clk(clk), .reset(n9), .execution_stage_out(alu_out), 
        .b_reg_out(b_reg_out_ex), .rd_reg_out(rd_out_ex) );
  MEMORY_STAGE_numbit32 MEMORY ( .alu_in(alu_out), .rd_reg_in(rd_out_ex), 
        .reset(n9), .clk(clk), .to_mem_stage_reg(to_mem_stage_reg), 
        .rd_reg_out(rd_out_mem), .memory_stage_out(memory_stage_out), 
        .alu_out(alu_out_mem) );
  WRITE_BACK_STAGE_N32 WRITEBACK ( .LMD(memory_stage_out), .ALUOUT(alu_out_mem), .RD_IN(rd_out_mem), .CONTROL(wb_control), .JAL_SEL(jal_sel), .RD_OUT(
        rd_out_wb), .WB_OUT(wb_stage_out) );
  BUF_X1 U1 ( .A(reset), .Z(n9) );
endmodule


module DLX ( clk, reset, npc_out_bpu, npc_out_if, instruction_fetched, ir_out, 
        rd_out_id, npc_out_id, a_reg_out, b_reg_out, imm_reg_out, alu_out, 
        rd_out_ex, b_reg_out_ex, rd_out_mem, memory_stage_out, alu_out_mem, 
        rd_out_wb, wb_stage_out, address_error, MUXA_CONTROL, MUXB_CONTROL, 
        ALU_OPCODE, DRAM_WE, DRAM_RE, WB_MUX_SEL, JAL_SEL, RF_WE, 
        alu_forwarding_one, mem_forwarding_one, alu_forwarding_two, 
        mem_forwarding_two, alu_forwarding_value, mem_forwarding_value );
  output [31:0] npc_out_bpu;
  output [31:0] npc_out_if;
  output [31:0] instruction_fetched;
  output [31:0] ir_out;
  output [4:0] rd_out_id;
  output [31:0] npc_out_id;
  output [31:0] a_reg_out;
  output [31:0] b_reg_out;
  output [31:0] imm_reg_out;
  output [31:0] alu_out;
  output [4:0] rd_out_ex;
  output [31:0] b_reg_out_ex;
  output [4:0] rd_out_mem;
  output [31:0] memory_stage_out;
  output [31:0] alu_out_mem;
  output [4:0] rd_out_wb;
  output [31:0] wb_stage_out;
  output [3:0] ALU_OPCODE;
  output [31:0] alu_forwarding_value;
  output [31:0] mem_forwarding_value;
  input clk, reset;
  output address_error, MUXA_CONTROL, MUXB_CONTROL, DRAM_WE, DRAM_RE,
         WB_MUX_SEL, JAL_SEL, RF_WE, alu_forwarding_one, mem_forwarding_one,
         alu_forwarding_two, mem_forwarding_two;

  assign MUXA_CONTROL = 1'b0;
  assign MUXB_CONTROL = 1'b0;
  assign ALU_OPCODE[3] = 1'b0;
  assign ALU_OPCODE[2] = 1'b0;
  assign ALU_OPCODE[1] = 1'b0;
  assign ALU_OPCODE[0] = 1'b0;
  assign DRAM_WE = 1'b0;
  assign DRAM_RE = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign JAL_SEL = 1'b0;
  assign RF_WE = 1'b0;

  CU_HARDWIRED CONTROL_I ( .OPCODE(ir_out[31:26]), .FUNC(ir_out[10:0]), .Clk(
        clk), .Rst(reset) );
  DATAPATH_numbit32 DATAPATH_I ( .clk(clk), .reset(reset), .write_enable(1'b0), 
        .mux_one_control(1'b0), .mux_two_control(1'b0), .alu_control({1'b0, 
        1'b0, 1'b0, 1'b0}), .to_ir({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .to_mem_stage_reg({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .wb_control(1'b0), .jal_sel(1'b0), .npc_out_if(npc_out_if), 
        .npc_out_bpu(npc_out_bpu), .instruction_fetched(instruction_fetched), 
        .ir_out(ir_out), .rd_out_id(rd_out_id), .npc_out_id(npc_out_id), 
        .a_reg_out(a_reg_out), .b_reg_out(b_reg_out), .imm_reg_out(imm_reg_out), .alu_out(alu_out), .rd_out_ex(rd_out_ex), .b_reg_out_ex(b_reg_out_ex), 
        .rd_out_mem(rd_out_mem), .memory_stage_out(memory_stage_out), 
        .alu_out_mem(alu_out_mem), .wb_stage_out(wb_stage_out), .rd_out_wb(
        rd_out_wb), .alu_forwarding_one(alu_forwarding_one), 
        .mem_forwarding_one(mem_forwarding_one), .alu_forwarding_two(
        alu_forwarding_two), .mem_forwarding_two(mem_forwarding_two), 
        .alu_forwarding_value(alu_forwarding_value), .mem_forwarding_value(
        mem_forwarding_value) );
endmodule

